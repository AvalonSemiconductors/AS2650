// This is the unpowered netlist.
module wrapped_as2650 (wb_clk_i,
    io_in,
    io_oeb,
    io_out,
    la_data_out);
 input wb_clk_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 output [63:0] la_data_out;

 wire net148;
 wire net153;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net149;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net150;
 wire net118;
 wire net119;
 wire net120;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net151;
 wire net152;
 wire net121;
 wire net126;
 wire net122;
 wire net123;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net124;
 wire net125;
 wire net159;
 wire net132;
 wire net160;
 wire net133;
 wire net161;
 wire net134;
 wire net162;
 wire net135;
 wire net163;
 wire net136;
 wire net164;
 wire net137;
 wire net165;
 wire net138;
 wire net166;
 wire net139;
 wire net140;
 wire net167;
 wire net141;
 wire net168;
 wire net142;
 wire net169;
 wire net143;
 wire net170;
 wire net144;
 wire net171;
 wire net145;
 wire net172;
 wire net146;
 wire net173;
 wire net147;
 wire net174;
 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire \as2650.addr_buff[0] ;
 wire \as2650.addr_buff[1] ;
 wire \as2650.addr_buff[2] ;
 wire \as2650.addr_buff[3] ;
 wire \as2650.addr_buff[4] ;
 wire \as2650.addr_buff[5] ;
 wire \as2650.addr_buff[6] ;
 wire \as2650.addr_buff[7] ;
 wire \as2650.alu_op[0] ;
 wire \as2650.alu_op[1] ;
 wire \as2650.alu_op[2] ;
 wire \as2650.cycle[0] ;
 wire \as2650.cycle[10] ;
 wire \as2650.cycle[11] ;
 wire \as2650.cycle[12] ;
 wire \as2650.cycle[13] ;
 wire \as2650.cycle[1] ;
 wire \as2650.cycle[2] ;
 wire \as2650.cycle[3] ;
 wire \as2650.cycle[4] ;
 wire \as2650.cycle[5] ;
 wire \as2650.cycle[6] ;
 wire \as2650.cycle[7] ;
 wire \as2650.cycle[8] ;
 wire \as2650.cycle[9] ;
 wire \as2650.holding_reg[0] ;
 wire \as2650.holding_reg[1] ;
 wire \as2650.holding_reg[2] ;
 wire \as2650.holding_reg[3] ;
 wire \as2650.holding_reg[4] ;
 wire \as2650.holding_reg[5] ;
 wire \as2650.holding_reg[6] ;
 wire \as2650.holding_reg[7] ;
 wire \as2650.idx_ctrl[0] ;
 wire \as2650.idx_ctrl[1] ;
 wire \as2650.ins_reg[0] ;
 wire \as2650.ins_reg[1] ;
 wire \as2650.ins_reg[2] ;
 wire \as2650.ins_reg[3] ;
 wire \as2650.ins_reg[4] ;
 wire \as2650.ivec[0] ;
 wire \as2650.ivec[1] ;
 wire \as2650.ivec[2] ;
 wire \as2650.ivec[3] ;
 wire \as2650.ivec[4] ;
 wire \as2650.ivec[5] ;
 wire \as2650.ivec[6] ;
 wire \as2650.ivec[7] ;
 wire \as2650.last_intr ;
 wire \as2650.prefixed ;
 wire \as2650.r0[0] ;
 wire \as2650.r0[1] ;
 wire \as2650.r0[2] ;
 wire \as2650.r0[3] ;
 wire \as2650.r0[4] ;
 wire \as2650.r0[5] ;
 wire \as2650.r0[6] ;
 wire \as2650.r0[7] ;
 wire \as2650.r123[0][0] ;
 wire \as2650.r123[0][1] ;
 wire \as2650.r123[0][2] ;
 wire \as2650.r123[0][3] ;
 wire \as2650.r123[0][4] ;
 wire \as2650.r123[0][5] ;
 wire \as2650.r123[0][6] ;
 wire \as2650.r123[0][7] ;
 wire \as2650.r123[1][0] ;
 wire \as2650.r123[1][1] ;
 wire \as2650.r123[1][2] ;
 wire \as2650.r123[1][3] ;
 wire \as2650.r123[1][4] ;
 wire \as2650.r123[1][5] ;
 wire \as2650.r123[1][6] ;
 wire \as2650.r123[1][7] ;
 wire \as2650.r123[2][0] ;
 wire \as2650.r123[2][1] ;
 wire \as2650.r123[2][2] ;
 wire \as2650.r123[2][3] ;
 wire \as2650.r123[2][4] ;
 wire \as2650.r123[2][5] ;
 wire \as2650.r123[2][6] ;
 wire \as2650.r123[2][7] ;
 wire \as2650.r123[3][0] ;
 wire \as2650.r123[3][1] ;
 wire \as2650.r123[3][2] ;
 wire \as2650.r123[3][3] ;
 wire \as2650.r123[3][4] ;
 wire \as2650.r123[3][5] ;
 wire \as2650.r123[3][6] ;
 wire \as2650.r123[3][7] ;
 wire \as2650.r123_2[0][0] ;
 wire \as2650.r123_2[0][1] ;
 wire \as2650.r123_2[0][2] ;
 wire \as2650.r123_2[0][3] ;
 wire \as2650.r123_2[0][4] ;
 wire \as2650.r123_2[0][5] ;
 wire \as2650.r123_2[0][6] ;
 wire \as2650.r123_2[0][7] ;
 wire \as2650.r123_2[1][0] ;
 wire \as2650.r123_2[1][1] ;
 wire \as2650.r123_2[1][2] ;
 wire \as2650.r123_2[1][3] ;
 wire \as2650.r123_2[1][4] ;
 wire \as2650.r123_2[1][5] ;
 wire \as2650.r123_2[1][6] ;
 wire \as2650.r123_2[1][7] ;
 wire \as2650.r123_2[2][0] ;
 wire \as2650.r123_2[2][1] ;
 wire \as2650.r123_2[2][2] ;
 wire \as2650.r123_2[2][3] ;
 wire \as2650.r123_2[2][4] ;
 wire \as2650.r123_2[2][5] ;
 wire \as2650.r123_2[2][6] ;
 wire \as2650.r123_2[2][7] ;
 wire \as2650.r123_2[3][0] ;
 wire \as2650.r123_2[3][1] ;
 wire \as2650.r123_2[3][2] ;
 wire \as2650.r123_2[3][3] ;
 wire \as2650.r123_2[3][4] ;
 wire \as2650.r123_2[3][5] ;
 wire \as2650.r123_2[3][6] ;
 wire \as2650.r123_2[3][7] ;
 wire \as2650.stack[0][0] ;
 wire \as2650.stack[0][10] ;
 wire \as2650.stack[0][11] ;
 wire \as2650.stack[0][12] ;
 wire \as2650.stack[0][13] ;
 wire \as2650.stack[0][14] ;
 wire \as2650.stack[0][1] ;
 wire \as2650.stack[0][2] ;
 wire \as2650.stack[0][3] ;
 wire \as2650.stack[0][4] ;
 wire \as2650.stack[0][5] ;
 wire \as2650.stack[0][6] ;
 wire \as2650.stack[0][7] ;
 wire \as2650.stack[0][8] ;
 wire \as2650.stack[0][9] ;
 wire \as2650.stack[10][0] ;
 wire \as2650.stack[10][10] ;
 wire \as2650.stack[10][11] ;
 wire \as2650.stack[10][12] ;
 wire \as2650.stack[10][13] ;
 wire \as2650.stack[10][14] ;
 wire \as2650.stack[10][1] ;
 wire \as2650.stack[10][2] ;
 wire \as2650.stack[10][3] ;
 wire \as2650.stack[10][4] ;
 wire \as2650.stack[10][5] ;
 wire \as2650.stack[10][6] ;
 wire \as2650.stack[10][7] ;
 wire \as2650.stack[10][8] ;
 wire \as2650.stack[10][9] ;
 wire \as2650.stack[11][0] ;
 wire \as2650.stack[11][10] ;
 wire \as2650.stack[11][11] ;
 wire \as2650.stack[11][12] ;
 wire \as2650.stack[11][13] ;
 wire \as2650.stack[11][14] ;
 wire \as2650.stack[11][1] ;
 wire \as2650.stack[11][2] ;
 wire \as2650.stack[11][3] ;
 wire \as2650.stack[11][4] ;
 wire \as2650.stack[11][5] ;
 wire \as2650.stack[11][6] ;
 wire \as2650.stack[11][7] ;
 wire \as2650.stack[11][8] ;
 wire \as2650.stack[11][9] ;
 wire \as2650.stack[12][0] ;
 wire \as2650.stack[12][10] ;
 wire \as2650.stack[12][11] ;
 wire \as2650.stack[12][12] ;
 wire \as2650.stack[12][13] ;
 wire \as2650.stack[12][14] ;
 wire \as2650.stack[12][1] ;
 wire \as2650.stack[12][2] ;
 wire \as2650.stack[12][3] ;
 wire \as2650.stack[12][4] ;
 wire \as2650.stack[12][5] ;
 wire \as2650.stack[12][6] ;
 wire \as2650.stack[12][7] ;
 wire \as2650.stack[12][8] ;
 wire \as2650.stack[12][9] ;
 wire \as2650.stack[13][0] ;
 wire \as2650.stack[13][10] ;
 wire \as2650.stack[13][11] ;
 wire \as2650.stack[13][12] ;
 wire \as2650.stack[13][13] ;
 wire \as2650.stack[13][14] ;
 wire \as2650.stack[13][1] ;
 wire \as2650.stack[13][2] ;
 wire \as2650.stack[13][3] ;
 wire \as2650.stack[13][4] ;
 wire \as2650.stack[13][5] ;
 wire \as2650.stack[13][6] ;
 wire \as2650.stack[13][7] ;
 wire \as2650.stack[13][8] ;
 wire \as2650.stack[13][9] ;
 wire \as2650.stack[14][0] ;
 wire \as2650.stack[14][10] ;
 wire \as2650.stack[14][11] ;
 wire \as2650.stack[14][12] ;
 wire \as2650.stack[14][13] ;
 wire \as2650.stack[14][14] ;
 wire \as2650.stack[14][1] ;
 wire \as2650.stack[14][2] ;
 wire \as2650.stack[14][3] ;
 wire \as2650.stack[14][4] ;
 wire \as2650.stack[14][5] ;
 wire \as2650.stack[14][6] ;
 wire \as2650.stack[14][7] ;
 wire \as2650.stack[14][8] ;
 wire \as2650.stack[14][9] ;
 wire \as2650.stack[15][0] ;
 wire \as2650.stack[15][10] ;
 wire \as2650.stack[15][11] ;
 wire \as2650.stack[15][12] ;
 wire \as2650.stack[15][13] ;
 wire \as2650.stack[15][14] ;
 wire \as2650.stack[15][1] ;
 wire \as2650.stack[15][2] ;
 wire \as2650.stack[15][3] ;
 wire \as2650.stack[15][4] ;
 wire \as2650.stack[15][5] ;
 wire \as2650.stack[15][6] ;
 wire \as2650.stack[15][7] ;
 wire \as2650.stack[15][8] ;
 wire \as2650.stack[15][9] ;
 wire \as2650.stack[1][0] ;
 wire \as2650.stack[1][10] ;
 wire \as2650.stack[1][11] ;
 wire \as2650.stack[1][12] ;
 wire \as2650.stack[1][13] ;
 wire \as2650.stack[1][14] ;
 wire \as2650.stack[1][1] ;
 wire \as2650.stack[1][2] ;
 wire \as2650.stack[1][3] ;
 wire \as2650.stack[1][4] ;
 wire \as2650.stack[1][5] ;
 wire \as2650.stack[1][6] ;
 wire \as2650.stack[1][7] ;
 wire \as2650.stack[1][8] ;
 wire \as2650.stack[1][9] ;
 wire \as2650.stack[2][0] ;
 wire \as2650.stack[2][10] ;
 wire \as2650.stack[2][11] ;
 wire \as2650.stack[2][12] ;
 wire \as2650.stack[2][13] ;
 wire \as2650.stack[2][14] ;
 wire \as2650.stack[2][1] ;
 wire \as2650.stack[2][2] ;
 wire \as2650.stack[2][3] ;
 wire \as2650.stack[2][4] ;
 wire \as2650.stack[2][5] ;
 wire \as2650.stack[2][6] ;
 wire \as2650.stack[2][7] ;
 wire \as2650.stack[2][8] ;
 wire \as2650.stack[2][9] ;
 wire \as2650.stack[3][0] ;
 wire \as2650.stack[3][10] ;
 wire \as2650.stack[3][11] ;
 wire \as2650.stack[3][12] ;
 wire \as2650.stack[3][13] ;
 wire \as2650.stack[3][14] ;
 wire \as2650.stack[3][1] ;
 wire \as2650.stack[3][2] ;
 wire \as2650.stack[3][3] ;
 wire \as2650.stack[3][4] ;
 wire \as2650.stack[3][5] ;
 wire \as2650.stack[3][6] ;
 wire \as2650.stack[3][7] ;
 wire \as2650.stack[3][8] ;
 wire \as2650.stack[3][9] ;
 wire \as2650.stack[4][0] ;
 wire \as2650.stack[4][10] ;
 wire \as2650.stack[4][11] ;
 wire \as2650.stack[4][12] ;
 wire \as2650.stack[4][13] ;
 wire \as2650.stack[4][14] ;
 wire \as2650.stack[4][1] ;
 wire \as2650.stack[4][2] ;
 wire \as2650.stack[4][3] ;
 wire \as2650.stack[4][4] ;
 wire \as2650.stack[4][5] ;
 wire \as2650.stack[4][6] ;
 wire \as2650.stack[4][7] ;
 wire \as2650.stack[4][8] ;
 wire \as2650.stack[4][9] ;
 wire \as2650.stack[5][0] ;
 wire \as2650.stack[5][10] ;
 wire \as2650.stack[5][11] ;
 wire \as2650.stack[5][12] ;
 wire \as2650.stack[5][13] ;
 wire \as2650.stack[5][14] ;
 wire \as2650.stack[5][1] ;
 wire \as2650.stack[5][2] ;
 wire \as2650.stack[5][3] ;
 wire \as2650.stack[5][4] ;
 wire \as2650.stack[5][5] ;
 wire \as2650.stack[5][6] ;
 wire \as2650.stack[5][7] ;
 wire \as2650.stack[5][8] ;
 wire \as2650.stack[5][9] ;
 wire \as2650.stack[6][0] ;
 wire \as2650.stack[6][10] ;
 wire \as2650.stack[6][11] ;
 wire \as2650.stack[6][12] ;
 wire \as2650.stack[6][13] ;
 wire \as2650.stack[6][14] ;
 wire \as2650.stack[6][1] ;
 wire \as2650.stack[6][2] ;
 wire \as2650.stack[6][3] ;
 wire \as2650.stack[6][4] ;
 wire \as2650.stack[6][5] ;
 wire \as2650.stack[6][6] ;
 wire \as2650.stack[6][7] ;
 wire \as2650.stack[6][8] ;
 wire \as2650.stack[6][9] ;
 wire \as2650.stack[7][0] ;
 wire \as2650.stack[7][10] ;
 wire \as2650.stack[7][11] ;
 wire \as2650.stack[7][12] ;
 wire \as2650.stack[7][13] ;
 wire \as2650.stack[7][14] ;
 wire \as2650.stack[7][1] ;
 wire \as2650.stack[7][2] ;
 wire \as2650.stack[7][3] ;
 wire \as2650.stack[7][4] ;
 wire \as2650.stack[7][5] ;
 wire \as2650.stack[7][6] ;
 wire \as2650.stack[7][7] ;
 wire \as2650.stack[7][8] ;
 wire \as2650.stack[7][9] ;
 wire \as2650.stack[8][0] ;
 wire \as2650.stack[8][10] ;
 wire \as2650.stack[8][11] ;
 wire \as2650.stack[8][12] ;
 wire \as2650.stack[8][13] ;
 wire \as2650.stack[8][14] ;
 wire \as2650.stack[8][1] ;
 wire \as2650.stack[8][2] ;
 wire \as2650.stack[8][3] ;
 wire \as2650.stack[8][4] ;
 wire \as2650.stack[8][5] ;
 wire \as2650.stack[8][6] ;
 wire \as2650.stack[8][7] ;
 wire \as2650.stack[8][8] ;
 wire \as2650.stack[8][9] ;
 wire \as2650.stack[9][0] ;
 wire \as2650.stack[9][10] ;
 wire \as2650.stack[9][11] ;
 wire \as2650.stack[9][12] ;
 wire \as2650.stack[9][13] ;
 wire \as2650.stack[9][14] ;
 wire \as2650.stack[9][1] ;
 wire \as2650.stack[9][2] ;
 wire \as2650.stack[9][3] ;
 wire \as2650.stack[9][4] ;
 wire \as2650.stack[9][5] ;
 wire \as2650.stack[9][6] ;
 wire \as2650.stack[9][7] ;
 wire \as2650.stack[9][8] ;
 wire \as2650.stack[9][9] ;
 wire clknet_0_wb_clk_i;
 wire clknet_3_0_0_wb_clk_i;
 wire clknet_3_1_0_wb_clk_i;
 wire clknet_3_2_0_wb_clk_i;
 wire clknet_3_3_0_wb_clk_i;
 wire clknet_3_4_0_wb_clk_i;
 wire clknet_3_5_0_wb_clk_i;
 wire clknet_3_6_0_wb_clk_i;
 wire clknet_3_7_0_wb_clk_i;
 wire clknet_4_0__leaf_wb_clk_i;
 wire clknet_4_10__leaf_wb_clk_i;
 wire clknet_4_11__leaf_wb_clk_i;
 wire clknet_4_12__leaf_wb_clk_i;
 wire clknet_4_13__leaf_wb_clk_i;
 wire clknet_4_14__leaf_wb_clk_i;
 wire clknet_4_15__leaf_wb_clk_i;
 wire clknet_4_1__leaf_wb_clk_i;
 wire clknet_4_2__leaf_wb_clk_i;
 wire clknet_4_3__leaf_wb_clk_i;
 wire clknet_4_4__leaf_wb_clk_i;
 wire clknet_4_5__leaf_wb_clk_i;
 wire clknet_4_6__leaf_wb_clk_i;
 wire clknet_4_7__leaf_wb_clk_i;
 wire clknet_4_8__leaf_wb_clk_i;
 wire clknet_4_9__leaf_wb_clk_i;
 wire clknet_leaf_0_wb_clk_i;
 wire clknet_leaf_100_wb_clk_i;
 wire clknet_leaf_102_wb_clk_i;
 wire clknet_leaf_103_wb_clk_i;
 wire clknet_leaf_104_wb_clk_i;
 wire clknet_leaf_105_wb_clk_i;
 wire clknet_leaf_106_wb_clk_i;
 wire clknet_leaf_107_wb_clk_i;
 wire clknet_leaf_109_wb_clk_i;
 wire clknet_leaf_10_wb_clk_i;
 wire clknet_leaf_111_wb_clk_i;
 wire clknet_leaf_112_wb_clk_i;
 wire clknet_leaf_113_wb_clk_i;
 wire clknet_leaf_114_wb_clk_i;
 wire clknet_leaf_115_wb_clk_i;
 wire clknet_leaf_116_wb_clk_i;
 wire clknet_leaf_117_wb_clk_i;
 wire clknet_leaf_118_wb_clk_i;
 wire clknet_leaf_119_wb_clk_i;
 wire clknet_leaf_11_wb_clk_i;
 wire clknet_leaf_120_wb_clk_i;
 wire clknet_leaf_123_wb_clk_i;
 wire clknet_leaf_125_wb_clk_i;
 wire clknet_leaf_126_wb_clk_i;
 wire clknet_leaf_127_wb_clk_i;
 wire clknet_leaf_12_wb_clk_i;
 wire clknet_leaf_13_wb_clk_i;
 wire clknet_leaf_14_wb_clk_i;
 wire clknet_leaf_15_wb_clk_i;
 wire clknet_leaf_16_wb_clk_i;
 wire clknet_leaf_17_wb_clk_i;
 wire clknet_leaf_18_wb_clk_i;
 wire clknet_leaf_19_wb_clk_i;
 wire clknet_leaf_1_wb_clk_i;
 wire clknet_leaf_20_wb_clk_i;
 wire clknet_leaf_21_wb_clk_i;
 wire clknet_leaf_22_wb_clk_i;
 wire clknet_leaf_23_wb_clk_i;
 wire clknet_leaf_24_wb_clk_i;
 wire clknet_leaf_25_wb_clk_i;
 wire clknet_leaf_26_wb_clk_i;
 wire clknet_leaf_27_wb_clk_i;
 wire clknet_leaf_28_wb_clk_i;
 wire clknet_leaf_29_wb_clk_i;
 wire clknet_leaf_2_wb_clk_i;
 wire clknet_leaf_31_wb_clk_i;
 wire clknet_leaf_32_wb_clk_i;
 wire clknet_leaf_33_wb_clk_i;
 wire clknet_leaf_34_wb_clk_i;
 wire clknet_leaf_35_wb_clk_i;
 wire clknet_leaf_36_wb_clk_i;
 wire clknet_leaf_37_wb_clk_i;
 wire clknet_leaf_38_wb_clk_i;
 wire clknet_leaf_39_wb_clk_i;
 wire clknet_leaf_3_wb_clk_i;
 wire clknet_leaf_40_wb_clk_i;
 wire clknet_leaf_41_wb_clk_i;
 wire clknet_leaf_42_wb_clk_i;
 wire clknet_leaf_43_wb_clk_i;
 wire clknet_leaf_44_wb_clk_i;
 wire clknet_leaf_46_wb_clk_i;
 wire clknet_leaf_48_wb_clk_i;
 wire clknet_leaf_49_wb_clk_i;
 wire clknet_leaf_4_wb_clk_i;
 wire clknet_leaf_50_wb_clk_i;
 wire clknet_leaf_52_wb_clk_i;
 wire clknet_leaf_53_wb_clk_i;
 wire clknet_leaf_58_wb_clk_i;
 wire clknet_leaf_59_wb_clk_i;
 wire clknet_leaf_5_wb_clk_i;
 wire clknet_leaf_60_wb_clk_i;
 wire clknet_leaf_61_wb_clk_i;
 wire clknet_leaf_63_wb_clk_i;
 wire clknet_leaf_64_wb_clk_i;
 wire clknet_leaf_65_wb_clk_i;
 wire clknet_leaf_66_wb_clk_i;
 wire clknet_leaf_67_wb_clk_i;
 wire clknet_leaf_68_wb_clk_i;
 wire clknet_leaf_69_wb_clk_i;
 wire clknet_leaf_6_wb_clk_i;
 wire clknet_leaf_70_wb_clk_i;
 wire clknet_leaf_71_wb_clk_i;
 wire clknet_leaf_72_wb_clk_i;
 wire clknet_leaf_73_wb_clk_i;
 wire clknet_leaf_74_wb_clk_i;
 wire clknet_leaf_75_wb_clk_i;
 wire clknet_leaf_76_wb_clk_i;
 wire clknet_leaf_77_wb_clk_i;
 wire clknet_leaf_78_wb_clk_i;
 wire clknet_leaf_79_wb_clk_i;
 wire clknet_leaf_7_wb_clk_i;
 wire clknet_leaf_81_wb_clk_i;
 wire clknet_leaf_82_wb_clk_i;
 wire clknet_leaf_83_wb_clk_i;
 wire clknet_leaf_84_wb_clk_i;
 wire clknet_leaf_85_wb_clk_i;
 wire clknet_leaf_86_wb_clk_i;
 wire clknet_leaf_87_wb_clk_i;
 wire clknet_leaf_8_wb_clk_i;
 wire clknet_leaf_91_wb_clk_i;
 wire clknet_leaf_92_wb_clk_i;
 wire clknet_leaf_93_wb_clk_i;
 wire clknet_leaf_94_wb_clk_i;
 wire clknet_leaf_95_wb_clk_i;
 wire clknet_leaf_96_wb_clk_i;
 wire clknet_leaf_97_wb_clk_i;
 wire clknet_leaf_98_wb_clk_i;
 wire clknet_leaf_99_wb_clk_i;
 wire clknet_leaf_9_wb_clk_i;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_1 (.I(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05862__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05863__I (.I(_05716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05865__I (.I(_05718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05866__I (.I(\as2650.ins_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05868__I (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05869__I (.I(\as2650.ins_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05870__I (.I(_05723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05872__A2 (.I(_05725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05873__I (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05874__I (.I(_05723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05875__A1 (.I(_05727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05875__A2 (.I(_05728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05876__I (.I(\as2650.ins_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05877__I (.I(_05730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05879__I (.I(_05732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05880__A1 (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05881__I (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05882__I (.I(_05732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05883__A1 (.I(_05735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05883__A2 (.I(_05736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05885__I (.I(\as2650.alu_op[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05887__I (.I(\as2650.alu_op[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05890__I (.I(_05743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05891__A1 (.I(_05728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05891__A2 (.I(_05736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05892__A1 (.I(_05745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05892__A2 (.I(_05738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05893__I (.I(\as2650.ins_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05895__A1 (.I(_05747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05896__A2 (.I(_05738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05896__A3 (.I(_05744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05896__B2 (.I(_05749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05897__I (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05898__I (.I(\as2650.ins_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05900__I (.I(_05753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05903__I (.I(\as2650.r0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05905__A1 (.I(_05723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05905__A2 (.I(_05730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05909__A1 (.I(_05728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05910__I (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05912__I (.I(_05765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05914__A1 (.I(_05758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05914__B1 (.I(_05763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05914__B2 (.I(_05767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05915__A1 (.I(\as2650.ins_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05915__A2 (.I(_05730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05920__I (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05923__I (.I(_05776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05925__A1 (.I(_05773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05925__A2 (.I(_05778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05927__I (.I(_05780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05928__A2 (.I(_05736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05929__A1 (.I(_05780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05929__A2 (.I(\as2650.r123[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05930__A1 (.I(_05781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05930__A2 (.I(\as2650.r123_2[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05930__B (.I(_05782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05931__A1 (.I(_05768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05932__I (.I(\as2650.r0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05933__I (.I(_05786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05934__A1 (.I(_05787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05935__S (.I(_05776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05936__I2 (.I(\as2650.r123_2[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05936__S1 (.I(_05776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05937__A1 (.I(\as2650.ins_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05937__A2 (.I(\as2650.ins_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05940__A2 (.I(_05789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05940__B1 (.I(_05790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05942__I (.I(\as2650.r0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05944__A1 (.I(_05797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05946__I (.I(_05799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05948__I1 (.I(\as2650.r123[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05948__I2 (.I(\as2650.r123_2[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05949__A2 (.I(_05801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05952__I (.I(\as2650.r0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05954__I (.I(_05807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05955__I (.I(_05808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05956__A1 (.I(_05809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05957__S (.I(_05776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05958__I1 (.I(\as2650.r123[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05958__I3 (.I(\as2650.r123_2[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05959__A2 (.I(_05811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05959__B1 (.I(_05812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05964__S0 (.I(_05730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05966__A1 (.I(_05817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05966__B2 (.I(_05818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05966__C1 (.I(_05819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05969__I (.I(\as2650.r0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05971__S0 (.I(\as2650.ins_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05973__A1 (.I(_05824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05973__B2 (.I(_05825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05973__C1 (.I(_05826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05975__A1 (.I(\as2650.ins_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05975__A2 (.I(\as2650.alu_op[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05975__A3 (.I(\as2650.alu_op[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05976__I (.I(\as2650.r0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05977__I3 (.I(\as2650.r123_2[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05977__S0 (.I(\as2650.ins_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05977__S1 (.I(_05799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05978__S (.I(_05799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05979__A1 (.I(_05830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05979__B2 (.I(_05831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05979__C1 (.I(_05832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05981__A2 (.I(_05829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05981__A3 (.I(_05834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05982__A3 (.I(_05835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05983__A1 (.I(_05805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05983__A2 (.I(_05814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05989__I (.I(_05842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05990__I (.I(_05829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05991__A2 (.I(_05844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05992__A1 (.I(_05841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05992__A2 (.I(_05845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05995__A1 (.I(_05809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05995__B2 (.I(_05812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05995__C1 (.I(_05811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05997__A2 (.I(_05850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05998__A2 (.I(_05851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__05999__A1 (.I(_05840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06000__I (.I(\as2650.r0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06001__I (.I(_05854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06002__A1 (.I(_05855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06004__I2 (.I(\as2650.r123_2[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06004__I3 (.I(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06004__S0 (.I(_05732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06006__A2 (.I(_05857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06008__S (.I(_05861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06009__A1 (.I(_05785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06012__A1 (.I(_00422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06013__I (.I(_05840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06014__A1 (.I(_00425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06020__A2 (.I(_00431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06021__A1 (.I(_05814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06022__I (.I(_05814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06023__A1 (.I(_00434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06024__A1 (.I(_00429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06026__I (.I(_05817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06027__A1 (.I(_00438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06028__A2 (.I(_05819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06028__B1 (.I(_05818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06030__I (.I(_00431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06031__I (.I(_05834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06033__I (.I(_00444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06034__A2 (.I(_00445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06034__A3 (.I(_05845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06036__A2 (.I(_05835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06037__A1 (.I(_00441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06039__A1 (.I(_05850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06041__A1 (.I(_05835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06043__A1 (.I(_05844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06043__A2 (.I(_00445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06044__A1 (.I(_00450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06044__A2 (.I(_00452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06044__A3 (.I(_00454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06044__A4 (.I(_00455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06045__A1 (.I(_00437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06046__A1 (.I(_00421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06046__A2 (.I(_00424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06046__A3 (.I(_00428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06047__A1 (.I(_05754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06047__A2 (.I(_05756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06047__A3 (.I(_00458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06048__A2 (.I(_00459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06052__I (.I(_00463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06053__A2 (.I(_05747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06055__I (.I(_00466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06058__I (.I(_00463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06060__A1 (.I(_05773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06060__A2 (.I(_00469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06061__I (.I(_00472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06062__A1 (.I(_05723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06062__A2 (.I(_05732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06065__A1 (.I(_00476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06066__A2 (.I(_00477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06068__I (.I(_00479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06070__A1 (.I(_00481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06070__A2 (.I(_00463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06071__A2 (.I(_00482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06072__A1 (.I(_00475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06072__A2 (.I(_00483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06073__I (.I(\as2650.prefixed ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06075__A1 (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06077__A2 (.I(_00488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06080__A1 (.I(_00473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06080__A2 (.I(_00491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06081__A2 (.I(_00462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06081__A3 (.I(_00467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06083__A1 (.I(_00494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06083__A3 (.I(_00482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06084__A1 (.I(_00495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06084__A2 (.I(_00488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06086__A1 (.I(_00496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06087__I (.I(_05716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06088__A1 (.I(_05842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06089__A1 (.I(_00479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06090__A2 (.I(_00501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06091__I (.I(_00502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06092__A2 (.I(_00503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06095__I (.I(_00506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06096__I (.I(_00479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06097__I (.I(_00508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06098__A1 (.I(_05745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06098__A2 (.I(_05743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06099__A1 (.I(_00509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06099__A2 (.I(_00510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06101__I (.I(_00512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06103__I (.I(_00488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06104__A1 (.I(\as2650.prefixed ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06105__A1 (.I(_00515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06105__A2 (.I(_00516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06107__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06109__I (.I(_05747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06110__A1 (.I(\as2650.prefixed ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06111__A2 (.I(_00522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06112__A2 (.I(_00523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06114__I (.I(_00481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06115__I (.I(_05842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06116__A1 (.I(_00526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06117__A1 (.I(_00525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06118__A2 (.I(_00529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06119__A1 (.I(_00507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06119__A2 (.I(_00514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06122__I (.I(_00533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06124__I (.I(_00535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06125__I (.I(_00536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06126__I (.I(_00537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06127__A2 (.I(_00505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06127__B (.I(_00538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06128__A1 (.I(_00508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06128__A2 (.I(_00472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06130__I (.I(_00541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06132__I (.I(_00516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06133__A1 (.I(_00515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06133__A2 (.I(_00544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06136__A1 (.I(_00543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06136__A2 (.I(_00547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06137__I (.I(\as2650.prefixed ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06138__A2 (.I(_05753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06142__A1 (.I(_00476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06143__A1 (.I(_05743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06144__A1 (.I(_00479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06144__A2 (.I(_00463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06145__I (.I(_00556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06149__A1 (.I(_00494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06149__A3 (.I(_00560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06150__A2 (.I(_05753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06151__A1 (.I(_00481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06151__A2 (.I(_05749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06153__A1 (.I(_00515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06153__A2 (.I(_00561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06156__A1 (.I(_00508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06157__A1 (.I(_00508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06157__A3 (.I(_05844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06158__A1 (.I(_00568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06159__A2 (.I(_00570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06160__A2 (.I(_00571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06161__A1 (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06164__I (.I(_00575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06165__A1 (.I(_00553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06165__B (.I(_00482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06165__C (.I(_00576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06169__I (.I(_00580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06172__I (.I(_00583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06173__A1 (.I(_00578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06173__A2 (.I(_00584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06175__A2 (.I(_00577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06178__I (.I(_00476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06180__A2 (.I(_00591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06181__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06183__A1 (.I(_00594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06185__I (.I(_00596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06186__I (.I(_00597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06188__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06191__I (.I(_00602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06192__I (.I(_00603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06193__A1 (.I(_00599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06193__A2 (.I(_00604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06194__A1 (.I(_00598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06198__I (.I(_00609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06200__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06204__I (.I(_00615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06205__A1 (.I(_00594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06208__A2 (.I(_00610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06211__A1 (.I(_00496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06211__A2 (.I(_00622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06213__I (.I(_05754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06214__I (.I(_00625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06215__I (.I(_00626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06216__I (.I(_00627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06217__I (.I(\as2650.addr_buff[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06218__I (.I(_00629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06219__I (.I(_00630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06220__I (.I(_00631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06224__I (.I(_00635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06227__A1 (.I(_00636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06227__A2 (.I(_00638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06228__A1 (.I(_00628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06228__A2 (.I(_00506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06229__A2 (.I(_00624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06229__B2 (.I(_00491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06231__A2 (.I(_00642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06236__A1 (.I(_00592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06236__A3 (.I(_00647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06238__A1 (.I(_00575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06239__A2 (.I(_00647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06240__A1 (.I(_00610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06240__A3 (.I(_00651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06244__A1 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06245__I (.I(_00656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06246__A2 (.I(_00657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06247__A1 (.I(_00472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06249__I (.I(_00660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06251__A1 (.I(_00594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06251__A2 (.I(_00662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06254__A1 (.I(_00654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06255__A1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06257__I (.I(_00522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06258__I (.I(_00568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06261__I (.I(_00656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06262__A2 (.I(_00673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06264__A2 (.I(_00675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06265__A1 (.I(_00671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06266__I (.I(_00509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06269__A1 (.I(_00678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06269__A2 (.I(_00679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06269__A3 (.I(_00680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06270__I (.I(_00681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06272__A1 (.I(_00678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06272__A2 (.I(_00683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06272__A3 (.I(_05844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06274__A2 (.I(_00685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06277__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06278__A3 (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06279__I (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06280__A1 (.I(_00688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06281__A1 (.I(_05716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06281__A2 (.I(_00692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06282__A1 (.I(_00668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06282__A2 (.I(_00677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06282__C (.I(_00693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06286__I (.I(_00697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06288__I (.I(_00657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06289__A1 (.I(_00512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06289__A2 (.I(_00700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06290__A1 (.I(_00594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06291__A2 (.I(_00701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06292__A1 (.I(_05716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06292__A2 (.I(_00699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06294__A3 (.I(_00681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06294__A4 (.I(_00570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06297__I (.I(_00708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06298__I (.I(_00709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06299__A1 (.I(_00695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06299__B2 (.I(_00710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06301__I (.I(_00642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06304__I (.I(_00510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06305__A1 (.I(_00526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06305__A2 (.I(_00715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06306__I (.I(_00716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06308__I (.I(_00718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06309__A1 (.I(_00719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06309__A2 (.I(_00491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06310__A1 (.I(\as2650.addr_buff[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06311__A2 (.I(_00467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06311__A4 (.I(_00721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06313__I (.I(_00723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06314__A1 (.I(_00679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06316__A1 (.I(_00724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06316__A2 (.I(_00726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06318__A2 (.I(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06320__A1 (.I(_00701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06320__A2 (.I(_00722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06322__A2 (.I(_00657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06323__I (.I(_00732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06324__I (.I(_00733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06325__I (.I(_00599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06327__A1 (.I(_00481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06327__A2 (.I(_00472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06329__I (.I(_00738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06331__I (.I(_00740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06332__I (.I(_00723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06334__A1 (.I(_00736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06334__A2 (.I(_00741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06334__A3 (.I(_00743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06335__A1 (.I(_00547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06335__A2 (.I(_00734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06336__I (.I(_00700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06339__I (.I(_00488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06340__A2 (.I(_00622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06341__A1 (.I(_00662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06341__A2 (.I(_00749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06342__A1 (.I(_00748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06343__B2 (.I(_00483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06346__I (.I(_00754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06347__A1 (.I(_00597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06352__A1 (.I(_00507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06353__B1 (.I(_00756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06356__I (.I(_00609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06357__I (.I(_00651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06362__A1 (.I(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06362__A3 (.I(_00769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06363__A1 (.I(_00736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06363__A2 (.I(_00766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06363__A3 (.I(_00770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06364__A1 (.I(_00764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06365__A2 (.I(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06366__I (.I(_00736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06368__I (.I(_00749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06371__A1 (.I(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06371__A2 (.I(_00777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06372__I (.I(\as2650.cycle[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06375__I (.I(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06376__I (.I(_00782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06378__A1 (.I(_00688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06379__A1 (.I(_00773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06380__I (.I(_00660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06382__A1 (.I(_00787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06382__A2 (.I(_00701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06383__A1 (.I(_00736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06383__A3 (.I(_00788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06384__B2 (.I(_00547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06386__I (.I(_00580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06387__I (.I(_00791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06388__I (.I(_00792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06389__I (.I(_00793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06390__I (.I(_00794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06391__I (.I(_00795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06396__A2 (.I(_00800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06398__A1 (.I(_00796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06398__A2 (.I(_00693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06398__B2 (.I(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06399__I (.I(_00803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06401__I (.I(_00804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06402__I (.I(_00805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06403__I (.I(_00622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06405__I (.I(_00808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06409__I (.I(_00812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06410__A1 (.I(_05754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06410__A2 (.I(_00477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06410__A3 (.I(_00813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06411__I (.I(_00814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06412__A1 (.I(_05842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06412__A2 (.I(_05747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06413__A1 (.I(_00680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06414__A2 (.I(_00807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06414__A3 (.I(_00815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06414__A4 (.I(_00817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06417__A1 (.I(_00494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06417__A2 (.I(_00820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06418__A2 (.I(_00591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06419__A1 (.I(_00525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06419__A2 (.I(_00822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06420__A1 (.I(_00813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06420__A2 (.I(_00823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06421__I (.I(_00626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06423__I (.I(_00826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06424__I (.I(_00678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06425__I (.I(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06426__I (.I(_00829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06427__I (.I(_00830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06429__I (.I(_00832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06431__A2 (.I(_00834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06433__I (.I(_00836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06434__I (.I(_00837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06435__I (.I(_00838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06436__I (.I(_00839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06437__A1 (.I(_00827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06437__C (.I(_00840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06438__B1 (.I(_00841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06438__B2 (.I(_00748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06439__A2 (.I(_00505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06440__A1 (.I(_00806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06440__A2 (.I(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06440__B1 (.I(_00842_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06440__B2 (.I(_00496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06441__I (.I(_00662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06442__I (.I(_00578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06443__I (.I(_00845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06444__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06446__I (.I(_00848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06447__I (.I(_00849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06448__I (.I(_00850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06449__I (.I(_00851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06451__I (.I(_00853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06454__I (.I(_00710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06455__I (.I(_00700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06456__A1 (.I(_00526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06457__I (.I(_00859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06458__I (.I(_00466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06459__A1 (.I(_00854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06459__A2 (.I(_00856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06459__B1 (.I(_00860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06459__B3 (.I(_00861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06460__A1 (.I(_00846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06460__A2 (.I(_00852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06460__A3 (.I(_00862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06461__A2 (.I(_00656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06462__I (.I(_00596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06464__A1 (.I(_05718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06464__B2 (.I(_00628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06465__A1 (.I(_00866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06466__A1 (.I(_00477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06467__A1 (.I(_00722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06467__A2 (.I(_00864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06468__A1 (.I(_00844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06468__A2 (.I(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06469__A2 (.I(_00807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06470__B1 (.I(_00871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06470__B2 (.I(_00576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06472__A1 (.I(_05754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06474__I (.I(_00874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06475__I (.I(_00875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06476__I (.I(_00876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06477__A2 (.I(_00877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06478__B1 (.I(_00873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06478__B2 (.I(_00878_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06481__A1 (.I(_00852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06481__A2 (.I(_00866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06482__I (.I(_00578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06484__A2 (.I(_00754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06485__A1 (.I(_00769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06485__A2 (.I(_00884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06486__A1 (.I(_00883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06486__A3 (.I(_00885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06488__A2 (.I(_00459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06490__A1 (.I(\as2650.addr_buff[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06490__A2 (.I(_00660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06491__A1 (.I(_00888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06491__A2 (.I(_00741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06491__B1 (.I(_00748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06491__B2 (.I(_00889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06492__A1 (.I(_00854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06492__A2 (.I(_00547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06493__I (.I(_00503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06494__I (.I(_00570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06496__I (.I(_00709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06497__A2 (.I(_00501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06499__A1 (.I(_00897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06500__A1 (.I(_00894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06500__A2 (.I(_00895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06501__A3 (.I(_00893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06502__I (.I(_00494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06504__I (.I(_00560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06505__A1 (.I(_00902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06509__A1 (.I(_00856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06509__A2 (.I(_00904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06509__A3 (.I(_00907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06511__A1 (.I(_00688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06511__A2 (.I(_00693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06511__C (.I(_00909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06512__A1 (.I(_00826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06512__A2 (.I(_00805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06512__A3 (.I(_00856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06512__B2 (.I(_00483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06515__I (.I(_00913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06518__I (.I(_00916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06521__A1 (.I(_00688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06521__A3 (.I(_00919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06524__A1 (.I(_00917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06525__A1 (.I(_00914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06525__A2 (.I(_00495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06525__B (.I(_00800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06525__C (.I(_00923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06528__I (.I(_00787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06530__A3 (.I(_00928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06530__A4 (.I(_00726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06531__A2 (.I(_00743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06531__A3 (.I(_00695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06534__A2 (.I(_00862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06535__A2 (.I(_00561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06536__A1 (.I(_00476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06536__A2 (.I(_05753_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06537__I (.I(_05782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06538__A1 (.I(_00936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06538__A2 (.I(_00560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06539__A2 (.I(_00937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06544__I (.I(_05744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06545__A1 (.I(_00943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06545__A3 (.I(_00937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06546__A1 (.I(_00939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06546__A2 (.I(_00942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06546__A3 (.I(_00944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06547__I (.I(_05773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06548__I (.I(_00946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06551__A1 (.I(_00947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06552__A1 (.I(_00624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06552__A2 (.I(_00823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06553__B (.I(_00950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06554__I (.I(_00522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06555__A1 (.I(_00575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06555__A2 (.I(_00953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06556__A1 (.I(_00680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06558__A3 (.I(_00954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06558__A4 (.I(_00956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06559__A2 (.I(_00815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06559__A3 (.I(_00956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06559__A4 (.I(_00904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06560__I (.I(_00953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06563__A1 (.I(_00678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06563__A3 (.I(_00961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06565__A2 (.I(_05749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06566__A1 (.I(_00946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06569__I (.I(_00967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06571__A1 (.I(_00800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06571__A2 (.I(_00963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06571__B1 (.I(_00965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06571__B2 (.I(_00969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06572__I (.I(_05736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06573__I (.I(_05728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06574__A2 (.I(_00812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06576__A2 (.I(_00974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06577__A2 (.I(_00975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06578__A1 (.I(_00960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06579__I (.I(_00561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06580__A1 (.I(_00837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06580__A2 (.I(_00978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06581__I (.I(_00820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06582__A1 (.I(_05763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06583__I (.I(_00981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06584__I (.I(_00982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06586__A1 (.I(_00856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06586__A2 (.I(_00984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06587__B2 (.I(_00668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06588__A1 (.I(_00496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06589__B (.I(_00538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06591__I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06592__I (.I(_00936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06593__A1 (.I(_05781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06593__A2 (.I(_00475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06595__A1 (.I(\as2650.cycle[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06595__A2 (.I(_00991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06597__A1 (.I(_00990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06597__A2 (.I(_00993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06599__A2 (.I(_00995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06600__I (.I(_05756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06601__A2 (.I(_00544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06602__A1 (.I(_00996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06603__A1 (.I(_05780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06604__A1 (.I(\as2650.cycle[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06605__I (.I(_01001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06606__A1 (.I(_00991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06606__A2 (.I(_00522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06607__A2 (.I(_01003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06608__A1 (.I(_00673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06608__A4 (.I(_01004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06610__I (.I(_05780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06611__I (.I(_01007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06614__A2 (.I(_01010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06617__A1 (.I(_00804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06617__A3 (.I(_01012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06617__A4 (.I(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06619__I (.I(_00991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06621__I (.I(_01017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06622__A1 (.I(_01008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06622__A2 (.I(_01014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06622__A3 (.I(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06623__C (.I(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06625__A2 (.I(_00993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06626__A1 (.I(_00814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06626__A2 (.I(_01021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06626__A3 (.I(_01022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06628__I (.I(_01010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06630__A2 (.I(_00916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06631__A1 (.I(_00615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06631__A2 (.I(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06631__A3 (.I(_01017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06631__A4 (.I(_01027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06632__A2 (.I(_00884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06633__A1 (.I(_01021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06633__A2 (.I(_01028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06633__A3 (.I(_01029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06634__A1 (.I(_00580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06635__A1 (.I(_00885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06637__A1 (.I(_01033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06637__A2 (.I(_00662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06637__A3 (.I(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06640__A1 (.I(_01035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06640__A2 (.I(_01036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06641__A1 (.I(\as2650.addr_buff[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06643__A1 (.I(_00990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06643__A2 (.I(_01032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06647__I (.I(_01043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06648__A1 (.I(_00989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06650__I (.I(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06653__A3 (.I(_05841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06654__I (.I(_01050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06655__I (.I(_05830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06656__I (.I(_01052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06657__I (.I(_01053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06659__A1 (.I(_00885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06660__A1 (.I(_01021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06661__I (.I(_01057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06663__I (.I(_00993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06665__A2 (.I(_01061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06667__A1 (.I(_00990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06667__A3 (.I(_01063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06668__I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06669__I (.I(_05785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06670__I (.I(_01066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06671__A1 (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06671__A2 (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06673__A1 (.I(_01065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06673__A2 (.I(_01067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06673__B (.I(_01069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06676__I (.I(_01072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06677__A2 (.I(_00568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06681__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06682__I (.I(_01078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06683__I (.I(_01079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06684__A1 (.I(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06685__A1 (.I(_00455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06690__A1 (.I(_01054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06691__A1 (.I(_00629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06692__A1 (.I(_00990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06692__A2 (.I(_01027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06692__A3 (.I(_01088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06692__A4 (.I(_01032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06696__A1 (.I(_05841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06697__I (.I(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06698__A2 (.I(_01094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06701__I0 (.I(_01051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06703__A1 (.I(_00445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06704__A1 (.I(_05773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06704__A2 (.I(_05832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06704__B1 (.I(_05831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06707__A2 (.I(_01103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06707__B (.I(_01052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06708__I (.I(_00808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06709__A1 (.I(_01101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06709__A2 (.I(_01103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06712__A1 (.I(_01108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06713__I (.I(_00683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06714__A3 (.I(_05756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06718__A1 (.I(_00444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06720__I (.I(_05744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06722__A1 (.I(_00683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06722__A3 (.I(_01118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06723__A1 (.I(_01117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06723__A2 (.I(_00961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06725__A2 (.I(_01109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06725__C (.I(_01121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06729__A2 (.I(_00943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06730__I (.I(_01126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06731__A1 (.I(_01069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06731__B (.I(_01127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06732__A1 (.I(_01069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06735__I (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06736__A1 (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06737__A2 (.I(_01133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06739__A2 (.I(_01133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06739__B (.I(_01135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06742__B2 (.I(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06743__A2 (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06744__A2 (.I(_01098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06745__I (.I(_01054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06746__I1 (.I(\as2650.r123_2[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06750__I (.I(_05781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06751__I (.I(_01022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06752__A1 (.I(_01147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06752__A2 (.I(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06753__A1 (.I(_00978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06754__I (.I(_01150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06755__A1 (.I(_01142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06755__A2 (.I(_01146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06756__A1 (.I(_00989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06756__C (.I(_00506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06759__A2 (.I(_01141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06761__I (.I(_01135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06762__B (.I(_01133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06763__A2 (.I(_00808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06764__A1 (.I(_00431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06766__A2 (.I(_05826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06766__B1 (.I(_05825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06768__I (.I(_05824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06769__A1 (.I(_01164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06769__B (.I(_00556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06770__A2 (.I(_00556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06770__B1 (.I(_01163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06783__A1 (.I(_01157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06784__I (.I(_00525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06785__A1 (.I(_01180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06785__A2 (.I(_00591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06786__A1 (.I(_01181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06787__C (.I(_01121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06790__B (.I(_01126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06792__B2 (.I(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06800__A1 (.I(_05841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06801__A1 (.I(_01192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06801__A2 (.I(_01196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06802__A1 (.I(_01192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06802__A2 (.I(_01196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06806__A1 (.I(_01035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06808__A1 (.I(_01192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06808__A2 (.I(_01203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06809__A1 (.I(_01192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06809__A2 (.I(_01203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06811__A2 (.I(_01206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06812__I (.I(_01164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06813__I (.I(_01208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06814__A1 (.I(_00815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06814__A2 (.I(_01021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06814__A3 (.I(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06816__I (.I(_01211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06817__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06819__I (.I(_01214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06820__I (.I(_01215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06821__A1 (.I(_00656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06821__A3 (.I(_01001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06821__A4 (.I(_01004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06823__A1 (.I(_00454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06824__A1 (.I(_01216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06827__A1 (.I(_01212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06828__I (.I(_00445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06829__I (.I(_01224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06830__A1 (.I(_01225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06831__A1 (.I(_01209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06833__A2 (.I(_01199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06834__I (.I(_01008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06836__A1 (.I(_01230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06836__A2 (.I(_01014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06836__A3 (.I(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06836__A4 (.I(_01231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06837__I0 (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06837__S (.I(_01232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06842__A1 (.I(_01053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06842__A2 (.I(_01237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06843__A1 (.I(_01208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06847__A2 (.I(_01233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06851__A1 (.I(_00431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06851__A2 (.I(_00444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06855__A3 (.I(_05834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06857__A2 (.I(_00444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06858__A2 (.I(_01251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06858__A3 (.I(_01252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06860__A1 (.I(_01251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06860__A2 (.I(_01252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06860__B (.I(_01035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06865__A2 (.I(_01259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06866__I (.I(_05850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06867__I (.I(_01261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06869__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06870__I (.I(_01264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06872__A1 (.I(_00450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06873__A1 (.I(_01265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06874__A1 (.I(_01262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06876__I (.I(_00438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06877__I (.I(_01271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06878__A1 (.I(_01272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06878__B (.I(_01057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06880__A2 (.I(_01260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06881__I0 (.I(_01254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06882__A2 (.I(_00525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06882__A3 (.I(_01118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06885__A1 (.I(_01211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06888__A2 (.I(_01010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06888__B2 (.I(_01271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06901__A1 (.I(_01277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06904__A1 (.I(_01109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06904__C (.I(_01121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06907__B (.I(_01127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06909__B2 (.I(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06910__I0 (.I(_01276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06910__I1 (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06910__S (.I(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06912__A1 (.I(_00438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06913__A1 (.I(_01164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06913__A2 (.I(_01237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06916__I (.I(_01310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06919__A1 (.I(_01052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06919__A2 (.I(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06925__A2 (.I(_01305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06926__A1 (.I(_05814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06928__A2 (.I(_01036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06929__A1 (.I(_05850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06929__B1 (.I(_01320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06930__I (.I(_05809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06931__I (.I(_01324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06933__I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06935__A1 (.I(_00452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06936__A1 (.I(_01328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06937__A1 (.I(_05805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06938__A1 (.I(_01211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06939__A1 (.I(_01325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06941__A2 (.I(_01323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06944__A1 (.I(_00434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06948__A2 (.I(_01320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06950__A2 (.I(_01343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06954__A1 (.I(_01261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06958__A2 (.I(_01010_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06958__B2 (.I(_01324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06967__A1 (.I(_01350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06967__A2 (.I(_01117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06968__I (.I(_01277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06975__B (.I(_01368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06976__A1 (.I(_00943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06976__A2 (.I(_00961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06977__A1 (.I(_01181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06980__A2 (.I(_01373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06985__A1 (.I(_05807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06989__I (.I(\as2650.r0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06990__I0 (.I(\as2650.r123[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06990__I1 (.I(\as2650.r123_2[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06990__S (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06991__I (.I(_01384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06992__I (.I(_01310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06993__A2 (.I(\as2650.r0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06995__I (.I(_01384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06998__A1 (.I(_05830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06998__A2 (.I(_01391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06998__B1 (.I(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__06998__B2 (.I(_05824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07005__A1 (.I(_05744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07006__I (.I(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07007__A1 (.I(_01147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07007__A2 (.I(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07008__I (.I(_01401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07011__A2 (.I(_01375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07011__B1 (.I(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07015__A4 (.I(_05834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07020__I (.I(_01412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07023__I (.I(_01415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07024__A2 (.I(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07025__I (.I(_05797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07027__I (.I(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07028__I (.I(_01420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07029__I (.I(_00425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07030__I (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07033__I (.I(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07034__A1 (.I(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07035__A1 (.I(_00437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07037__A1 (.I(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07038__A1 (.I(_01262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07039__A1 (.I(_01421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07041__A2 (.I(_01413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07043__A1 (.I(_00429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07045__A1 (.I(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07045__B1 (.I(_01012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07045__B2 (.I(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07054__A1 (.I(_01127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07061__A1 (.I(_01157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07064__A1 (.I(_01368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07064__B2 (.I(_01109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07069__I1 (.I(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07069__S (.I(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07074__I0 (.I(\as2650.r123[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07074__S (.I(_05799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07075__I (.I(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07076__A1 (.I(_01052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07080__A1 (.I(\as2650.r0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07081__A1 (.I(\as2650.r0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07084__A1 (.I(_05824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07094__A2 (.I(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07094__B1 (.I(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07095__I (.I(_01232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07096__A1 (.I(_00425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07101__I (.I(_05787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07102__B1 (.I(_01012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07105__A2 (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07107__I (.I(_00429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07108__A1 (.I(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07108__A2 (.I(_00812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07113__I (.I(_01127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07116__A2 (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07117__A2 (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07119__A1 (.I(_01181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07124__A1 (.I(_05840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07125__A1 (.I(_00429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07125__A2 (.I(_01261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07125__A3 (.I(_01251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07128__A1 (.I(_05805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07129__A1 (.I(_05840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07131__A1 (.I(_01522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07134__I (.I(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07138__A1 (.I(_01522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07139__I (.I(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07140__A2 (.I(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07142__I (.I(_00422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07143__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07144__I (.I(_01535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07145__A1 (.I(_00428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07146__A1 (.I(_01536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07147__A1 (.I(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07148__A1 (.I(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07149__A1 (.I(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07151__A2 (.I(_01526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07153__A2 (.I(_01514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07166__A1 (.I(_05830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07168__A1 (.I(_01164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07172__A1 (.I(\as2650.r0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07173__A1 (.I(_05786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07175__A1 (.I(\as2650.r0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07175__A4 (.I(_01310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07187__B1 (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07188__A2 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07189__I (.I(_05861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07192__A1 (.I(\as2650.holding_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07193__A1 (.I(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07196__I (.I(_05855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07197__B1 (.I(_01012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07198__A1 (.I(\as2650.holding_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07198__A2 (.I(_00820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07199__A1 (.I(_00820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07199__A2 (.I(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07204__A2 (.I(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07207__A1 (.I(_01157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07211__A1 (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07211__B (.I(_01350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07213__A1 (.I(_01109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07213__C (.I(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07216__A1 (.I(_00422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07219__A1 (.I(_05861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07219__A2 (.I(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07220__A2 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07221__A1 (.I(_00422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07223__I (.I(_01613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07225__I (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07226__I (.I(_01522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07227__A1 (.I(_05768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07228__A1 (.I(_00424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07229__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07232__I (.I(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07233__I (.I(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07234__A1 (.I(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07236__A1 (.I(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07237__A1 (.I(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07238__A1 (.I(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07238__B (.I(_01057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07239__C1 (.I(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07240__I (.I(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07241__A2 (.I(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07243__A2 (.I(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07244__A1 (.I(_01232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07245__A2 (.I(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07250__A1 (.I(_01208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07250__A2 (.I(_01640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07259__A1 (.I(_05817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07259__A2 (.I(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07263__I1 (.I(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07264__A1 (.I(\as2650.r0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07264__A2 (.I(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07265__A1 (.I(\as2650.r0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07266__A1 (.I(_05854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07268__A1 (.I(_05807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07268__A2 (.I(_01391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07278__B1 (.I(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07279__A2 (.I(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07281__A1 (.I(_01066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07283__I (.I(_05758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07285__A1 (.I(_01066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07285__A2 (.I(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07286__A1 (.I(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07286__A2 (.I(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07286__C (.I(_00812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07287__A2 (.I(_00560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07288__A1 (.I(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07290__A2 (.I(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07300__B (.I(_01368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07301__A1 (.I(_01181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07302__A1 (.I(_01121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07306__A1 (.I(_05785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07307__A2 (.I(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07308__A1 (.I(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07308__A2 (.I(_01697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07309__A1 (.I(_01066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07312__I (.I(_01701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07313__I (.I(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07314__A1 (.I(_01065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07314__A2 (.I(_01224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07314__B (.I(_01069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07316__A1 (.I(_00421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07317__A1 (.I(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07319__A1 (.I(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07320__A1 (.I(_01703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07320__B (.I(_01057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07322__A1 (.I(_01067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07323__I (.I(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07324__A2 (.I(_01713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07326__A2 (.I(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07327__A1 (.I(_01232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07328__A2 (.I(_01694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07334__I (.I(_01640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07335__A1 (.I(_00438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07335__A2 (.I(_01724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07344__A1 (.I(_05817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07344__A2 (.I(_01733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07346__A1 (.I(_05808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07346__A2 (.I(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07352__I (.I(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07354__A1 (.I(_05854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07357__A1 (.I(\as2650.r0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07357__A2 (.I(_01310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07358__A1 (.I(\as2650.r0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07358__A2 (.I(_01384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07359__A1 (.I(\as2650.r0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07359__A2 (.I(_05765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07369__A1 (.I(\as2650.r123[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07370__A2 (.I(_01718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07370__B1 (.I(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07372__I (.I(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07373__I (.I(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07374__I (.I(_01001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07376__A1 (.I(_00836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07376__A2 (.I(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07376__A3 (.I(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07377__I (.I(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07378__I (.I(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07379__I (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07381__I (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07382__A1 (.I(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07383__I (.I(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07384__I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07387__I (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07389__A1 (.I(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07390__I (.I(_01778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07394__I (.I(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07397__I (.I(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07399__A1 (.I(_01787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07399__A2 (.I(_01022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07400__A2 (.I(_01788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07401__A3 (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07402__A1 (.I(_00515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07403__A1 (.I(_00578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07403__A2 (.I(_01791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07405__A1 (.I(_00509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07405__A2 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07407__A1 (.I(_00889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07408__A1 (.I(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07408__B2 (.I(_00864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07409__A2 (.I(_00874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07410__A2 (.I(_05756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07411__A1 (.I(_01798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07411__A2 (.I(_01799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07412__A1 (.I(_00683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07414__A2 (.I(_00697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07415__B1 (.I(_01801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07416__A1 (.I(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07417__A1 (.I(_01789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07417__A2 (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07417__A3 (.I(_01805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07418__I (.I(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07419__I (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07421__I (.I(_01809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07423__I (.I(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07426__I (.I(_01814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07427__I (.I(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07428__A2 (.I(_01785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07429__I (.I(_01817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07430__A1 (.I(\as2650.stack[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07431__A1 (.I(_01789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07431__A2 (.I(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07431__A3 (.I(_01805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07432__I (.I(_01820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07433__I (.I(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07434__I (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07435__A1 (.I(_01822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07435__A2 (.I(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07436__I (.I(_01824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07438__I (.I(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07440__I (.I(_01053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07442__I (.I(_01789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07444__I (.I(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07445__I (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07446__I (.I(_01834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07449__A1 (.I(_01836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07450__A1 (.I(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07450__B (.I(_01838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07451__I (.I(_01839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07453__I (.I(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07454__A2 (.I(_01840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07455__A2 (.I(_01782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07455__B2 (.I(_01843_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07456__I (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07458__I (.I(_01845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07459__I (.I(_01846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07460__A1 (.I(\as2650.stack[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07461__I (.I(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07462__I (.I(_01209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07463__I (.I(_01850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07465__I (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07466__I (.I(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07468__A1 (.I(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07469__A1 (.I(_01851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07469__A2 (.I(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07470__I (.I(_01857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07471__I (.I(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07472__A1 (.I(_01849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07472__B (.I(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07473__A2 (.I(_01782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07474__I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07475__I (.I(_01861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07476__I (.I(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07478__I (.I(_01272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07479__I (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07480__I (.I(_01866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07482__I0 (.I(_01865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07482__I1 (.I(_01868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07482__S (.I(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07483__I (.I(_01869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07484__A1 (.I(_01849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07484__A2 (.I(_01870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07484__B (.I(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07485__A2 (.I(_01782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07486__I (.I(_01065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07487__I (.I(_01872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07488__I (.I(_01873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07489__A1 (.I(\as2650.stack[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07490__I (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07493__A1 (.I(_01325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07494__A1 (.I(_01877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07495__I (.I(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07496__A1 (.I(_01849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07496__A2 (.I(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07496__B (.I(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07497__A2 (.I(_01782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07498__I (.I(_01147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07499__I (.I(_01883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07500__I (.I(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07501__I (.I(_01817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07502__A1 (.I(\as2650.stack[13][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07503__I (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07505__A1 (.I(_01421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07505__A2 (.I(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07506__A1 (.I(_01889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07507__I (.I(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07508__A1 (.I(_01849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07508__A2 (.I(_01892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07508__B (.I(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07509__A1 (.I(_01884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07510__I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07512__I (.I(_01895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07514__I (.I(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07515__I (.I(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07516__I (.I(_01899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07517__I (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07518__I (.I(_01901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07520__A1 (.I(_01903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07521__A1 (.I(_01900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07521__A2 (.I(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07522__I (.I(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07523__A1 (.I(_01898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07524__A1 (.I(_01896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07525__I (.I(_05735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07526__I (.I(_01908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07527__A1 (.I(\as2650.stack[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07528__I (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07529__I (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07530__I (.I(_01912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07531__A1 (.I(_01913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07532__A1 (.I(_01911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07532__A2 (.I(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07532__B (.I(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07533__I (.I(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07534__A1 (.I(_01898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07535__A1 (.I(_01909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07536__I (.I(_05727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07537__I (.I(_01918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07539__I (.I(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07540__I (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07541__A1 (.I(_01922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07542__A1 (.I(_01921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07542__A2 (.I(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07542__B (.I(_01923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07543__I (.I(_01924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07544__A1 (.I(_01898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07545__A1 (.I(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07547__I (.I(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07548__I (.I(_01928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07549__I (.I(_01929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07550__A2 (.I(_00984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07551__A1 (.I(_01150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07553__A1 (.I(_01147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07553__A2 (.I(_00942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07555__I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07556__A1 (.I(_01936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07556__A2 (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07557__A1 (.I(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07558__A1 (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07558__A2 (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07560__A1 (.I(_01936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07560__B (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07562__I (.I(_01942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07563__I (.I(_01943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07564__I (.I(_01944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07565__A1 (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07569__I (.I(_01949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07572__I (.I(_01952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07573__I (.I(_01953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07574__I (.I(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07576__A2 (.I(_01951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07576__B1 (.I(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07576__B2 (.I(\as2650.stack[9][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07579__I (.I(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07580__I (.I(_01960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07584__I (.I(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07585__I (.I(_01965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07586__A2 (.I(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07586__B1 (.I(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07587__A1 (.I(_01950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07590__I (.I(_01970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07591__A2 (.I(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07591__B1 (.I(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07592__A2 (.I(_01951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07592__B1 (.I(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07593__A1 (.I(_01971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07597__A2 (.I(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07597__B1 (.I(_01977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07597__B2 (.I(\as2650.stack[1][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07600__I (.I(_01980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07601__I (.I(_01965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07602__A1 (.I(\as2650.stack[3][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07602__A2 (.I(_01981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07602__B2 (.I(\as2650.stack[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07603__A1 (.I(_01950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07604__I (.I(_01980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07605__B2 (.I(\as2650.stack[6][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07606__A1 (.I(\as2650.stack[4][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07606__A2 (.I(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07606__B1 (.I(_01977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07606__B2 (.I(\as2650.stack[5][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07607__A1 (.I(_01971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07609__A2 (.I(_01975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07610__A2 (.I(_01990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07613__A1 (.I(_01142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07614__A1 (.I(_05763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07614__A2 (.I(_01043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07616__B2 (.I(_01141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07617__A1 (.I(_05718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07620__I1 (.I(_01997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07623__I (.I(_01950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07624__I (.I(_01951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07625__I (.I(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07626__A2 (.I(_02004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07626__B1 (.I(_02005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07627__I (.I(_01981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07628__I (.I(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07629__A2 (.I(_02007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07629__B1 (.I(_02008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07630__A1 (.I(_02003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07631__I (.I(_01971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07632__I (.I(_01981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07634__A2 (.I(_02012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07634__B1 (.I(_02013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07635__I (.I(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07636__I (.I(_01977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07637__A2 (.I(_02015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07637__B1 (.I(_02016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07640__I (.I(_01949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07641__I (.I(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07642__I (.I(_01977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07643__A2 (.I(_02021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07643__B1 (.I(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07646__A2 (.I(_02024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07646__B1 (.I(_02025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07647__A1 (.I(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07648__I (.I(_01971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07652__I (.I(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07653__I (.I(_02032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07654__B1 (.I(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07658__B1 (.I(_02037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07659__A1 (.I(_02028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07659__A3 (.I(_02038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07660__I (.I(_01944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07661__B (.I(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07662__A2 (.I(_02019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07663__A2 (.I(_02042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07664__A1 (.I(_01850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07665__B2 (.I(_01233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07666__I1 (.I(_02045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07668__A2 (.I(_02004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07668__B1 (.I(_02005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07669__A2 (.I(_02007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07669__B1 (.I(_02008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07670__A1 (.I(_02003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07671__A2 (.I(_02012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07671__B1 (.I(_02013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07672__A2 (.I(_02015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07672__B1 (.I(_02016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07676__A2 (.I(_02054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07676__B1 (.I(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07677__I (.I(_02032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07678__A2 (.I(_02024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07679__A1 (.I(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07681__A2 (.I(_02059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07681__B1 (.I(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07683__B1 (.I(_02061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07684__A1 (.I(_02028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07684__A3 (.I(_02062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07685__B (.I(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07686__A2 (.I(_02053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07687__A2 (.I(_02065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07688__I (.I(_01272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07689__A1 (.I(_02067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07690__B2 (.I(_01305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07691__I1 (.I(_02069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07694__A2 (.I(_02021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07694__B1 (.I(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07695__A2 (.I(_02024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07695__B1 (.I(_02025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07696__A1 (.I(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07697__A2 (.I(_02024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07697__B1 (.I(_02025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07698__A2 (.I(_02021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07698__B1 (.I(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07701__I (.I(_01949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07703__A2 (.I(_01814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07703__B1 (.I(_02080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07703__B2 (.I(\as2650.stack[1][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07704__I (.I(_01960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07705__I (.I(_02032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07706__A2 (.I(_02082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07706__B1 (.I(_02083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07706__B2 (.I(\as2650.stack[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07708__I (.I(_01970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07709__I (.I(_01960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07710__A2 (.I(_02087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07710__B1 (.I(_02083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07713__A2 (.I(_02089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07713__B1 (.I(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07715__I (.I(_01944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07716__B (.I(_02093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07717__A2 (.I(_02078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07718__A2 (.I(_02095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07719__I (.I(_01325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07720__I (.I(_02097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07722__A1 (.I(_02098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07724__B2 (.I(_01375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07725__I0 (.I(\as2650.r123[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07725__I1 (.I(_02102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07727__A2 (.I(_02015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07727__B1 (.I(_02005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07728__A2 (.I(_02012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07728__B1 (.I(_02008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07729__A1 (.I(_02003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07729__A2 (.I(_02104_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07730__A2 (.I(_02012_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07730__B1 (.I(_02013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07731__A2 (.I(_02015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07731__B1 (.I(_02016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07734__A2 (.I(_02054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07734__B1 (.I(_02037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07736__A1 (.I(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07737__A2 (.I(_02059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07737__B1 (.I(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07738__B1 (.I(_02061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07739__A1 (.I(_02028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07740__B (.I(_02093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07742__A2 (.I(_02118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07743__I (.I(_01421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07744__A1 (.I(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07745__B2 (.I(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07747__I0 (.I(\as2650.r123[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07749__A1 (.I(\as2650.stack[8][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07749__A2 (.I(_02089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07749__B1 (.I(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07749__B2 (.I(\as2650.stack[9][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07750__I (.I(_02032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07751__A2 (.I(_02087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07751__B1 (.I(_02126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07753__I (.I(_01960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07754__A1 (.I(\as2650.stack[15][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07754__A2 (.I(_02129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07754__B1 (.I(_02126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07757__A1 (.I(\as2650.stack[12][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07757__A2 (.I(_02131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07757__B1 (.I(_02132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07760__A2 (.I(_02131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07760__B1 (.I(_02132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07761__I (.I(_01965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07762__A2 (.I(_02129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07762__B1 (.I(_02137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07762__B2 (.I(\as2650.stack[2][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07763__A1 (.I(_01950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07764__A2 (.I(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07764__B1 (.I(_02137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07765__A2 (.I(_01951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07765__B1 (.I(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07765__B2 (.I(\as2650.stack[5][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07768__A1 (.I(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07769__A2 (.I(_02144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07770__I (.I(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07771__A1 (.I(_02146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07772__B2 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07775__A2 (.I(_02054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07775__B1 (.I(_02037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07775__B2 (.I(\as2650.stack[9][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07779__A1 (.I(\as2650.stack[12][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07779__A2 (.I(_02054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07779__B1 (.I(_02037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07780__A1 (.I(_02028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07782__A2 (.I(_01814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07782__B1 (.I(_02080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07783__A2 (.I(_02082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07783__B1 (.I(_02083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07785__A2 (.I(_02087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07785__B1 (.I(_02126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07786__A2 (.I(_02089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07786__B1 (.I(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07786__B2 (.I(\as2650.stack[5][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07788__B (.I(_02093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07789__A1 (.I(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07790__A2 (.I(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07791__A1 (.I(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07792__B2 (.I(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07795__A1 (.I(_01921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07795__B1 (.I(_01718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07798__I (.I(_01820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07801__A2 (.I(_02173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07802__I (.I(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07804__I (.I(_02176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07806__I (.I(_01788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07808__I (.I(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07809__I (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07813__A1 (.I(_01146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07813__B2 (.I(_02185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07814__I (.I(_02186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07815__I (.I(_02176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07816__A2 (.I(_02188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07817__I (.I(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07818__I (.I(_01824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07819__A2 (.I(_01778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07819__A3 (.I(_02191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07821__I (.I(_02193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07823__I (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07825__I (.I(_02196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07826__A1 (.I(_01237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07826__B2 (.I(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07827__I (.I(_02198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07828__I (.I(_02176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07829__A2 (.I(_02200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07831__I (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07833__I (.I(_02203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07834__A1 (.I(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07834__B2 (.I(_02204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07835__I (.I(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07836__A2 (.I(_02200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07838__I (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07840__I (.I(_02209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07841__A1 (.I(_01391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07841__B2 (.I(_02210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07842__I (.I(_02211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07843__A2 (.I(_02200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07846__I (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07848__I (.I(_02216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07849__A1 (.I(_01724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07849__B2 (.I(_02217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07850__I (.I(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07851__A2 (.I(_02200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07852__I (.I(_02193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07854__I (.I(_01733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07856__I (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07857__A1 (.I(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07857__B2 (.I(_02224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07858__I (.I(_02225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07864__I (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07865__A1 (.I(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07865__B2 (.I(_02231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07866__I (.I(_02232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07870__A2 (.I(_01898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07871__I (.I(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07873__I (.I(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07887__I (.I(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07888__A2 (.I(_02191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07888__A3 (.I(_02246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07891__I (.I(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07893__A2 (.I(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07895__I (.I(_02080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07897__A1 (.I(_02250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07897__A2 (.I(_02253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07897__A3 (.I(_02255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07898__I (.I(_02256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07899__A1 (.I(\as2650.stack[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07900__I (.I(_01839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07902__A2 (.I(_02246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07903__I (.I(_02261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07906__I (.I(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07907__A1 (.I(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07908__A2 (.I(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07908__B2 (.I(_02266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07909__A1 (.I(\as2650.stack[10][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07910__I (.I(_01857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07911__I (.I(_02261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07912__I (.I(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07913__A1 (.I(_02268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07913__A2 (.I(_02269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07913__B (.I(_02270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07914__A2 (.I(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07915__A1 (.I(\as2650.stack[10][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07916__I (.I(_01869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07917__A1 (.I(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07917__A2 (.I(_02269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07917__B (.I(_02270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07918__A2 (.I(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07919__A1 (.I(\as2650.stack[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07920__I (.I(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07921__A1 (.I(_02276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07921__A2 (.I(_02269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07921__B (.I(_02270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07922__A2 (.I(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07923__I (.I(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07924__I (.I(_02256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07926__I (.I(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07927__A1 (.I(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07927__A2 (.I(_02269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07927__B (.I(_02270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07928__A1 (.I(_01884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07930__I (.I(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07931__I (.I(_02261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07932__A2 (.I(_02285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07933__A1 (.I(_01896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07934__A1 (.I(\as2650.stack[10][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07935__I (.I(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07936__A2 (.I(_02285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07937__A1 (.I(_01909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07939__I (.I(_01924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07940__A2 (.I(_02285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07941__A1 (.I(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07943__I (.I(_02293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07945__I (.I(_02293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07946__A2 (.I(_02296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07947__A2 (.I(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07948__I (.I(_02298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07949__A2 (.I(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07949__A3 (.I(_02299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07951__I (.I(_02301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07953__I (.I(_02293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07962__I (.I(_02301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07964__A1 (.I(\as2650.stack[12][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07966__A1 (.I(\as2650.stack[12][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07969__A2 (.I(_02246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07969__A3 (.I(_02299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07970__I (.I(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07971__I (.I(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07972__I (.I(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07973__A2 (.I(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07974__I (.I(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07975__A2 (.I(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07975__A3 (.I(_02318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07977__I (.I(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07979__I (.I(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07980__A2 (.I(_02322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07982__A2 (.I(_02322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07984__A2 (.I(_02322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07986__I (.I(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07987__A2 (.I(_02322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07988__I (.I(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07990__A2 (.I(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07992__A2 (.I(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07996__A1 (.I(_00836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07997__I (.I(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__07998__I (.I(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08000__A1 (.I(_00509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08000__A2 (.I(_00874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08001__A2 (.I(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08003__I (.I(_02339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08004__A1 (.I(_00584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08004__A2 (.I(_00944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08004__B1 (.I(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08006__A1 (.I(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08007__A1 (.I(_00936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08008__A1 (.I(_01703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08008__A2 (.I(_00535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08009__I (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08011__A1 (.I(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08011__A2 (.I(_00851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08012__A1 (.I(_00851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08013__A1 (.I(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08014__A2 (.I(_02345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08015__A1 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08015__A2 (.I(_02343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08015__B2 (.I(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08016__A1 (.I(_00773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08019__A2 (.I(_01785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08019__A4 (.I(_02255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08020__I (.I(_02355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08021__A1 (.I(\as2650.stack[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08022__A1 (.I(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08023__A2 (.I(_02354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08023__B2 (.I(_02358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08024__A1 (.I(\as2650.stack[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08025__I (.I(_02176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08026__I (.I(_02193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08027__A1 (.I(_02268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08027__A2 (.I(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08027__B (.I(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08028__A2 (.I(_02354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08030__A1 (.I(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08030__A2 (.I(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08030__B (.I(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08031__A2 (.I(_02354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08033__A1 (.I(_02276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08033__A2 (.I(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08033__B (.I(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08034__A2 (.I(_02354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08035__I (.I(_02193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08036__I (.I(_02355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08038__A1 (.I(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08038__A2 (.I(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08038__B (.I(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08039__A1 (.I(_01884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08041__A2 (.I(_02188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08042__A1 (.I(_01896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08043__A1 (.I(\as2650.stack[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08044__A2 (.I(_02188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08045__A1 (.I(_01909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08047__A2 (.I(_02188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08048__A1 (.I(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08049__I (.I(_02186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08051__A2 (.I(_02285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08052__I (.I(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08053__A1 (.I(_02377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08053__A2 (.I(_02378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08053__C (.I(_02380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08054__I (.I(_02198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08055__I (.I(_02261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08056__A2 (.I(_02382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08057__A1 (.I(_02381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08057__A2 (.I(_02378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08057__C (.I(_02380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08058__I (.I(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08059__A2 (.I(_02382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08060__A1 (.I(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08060__A2 (.I(_02378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08060__C (.I(_02380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08061__I (.I(_02211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08062__A2 (.I(_02382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08063__A1 (.I(_02386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08063__A2 (.I(_02378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08063__C (.I(_02380_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08064__I (.I(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08065__A2 (.I(_02382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08066__A1 (.I(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08067__I (.I(_02225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08069__A1 (.I(_02390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08070__I (.I(_02232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08072__A1 (.I(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08073__I (.I(_02137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08075__A2 (.I(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08078__I (.I(_02007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08079__I (.I(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08080__A1 (.I(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08082__A1 (.I(_02399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08083__I (.I(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08084__A1 (.I(\as2650.stack[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08085__I (.I(_01936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08086__A1 (.I(_02406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08086__A2 (.I(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08087__I (.I(_02407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08089__I (.I(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08092__I (.I(_02412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08093__A1 (.I(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08094__A2 (.I(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08094__B2 (.I(_02414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08096__I (.I(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08097__I (.I(_02412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08098__A1 (.I(_02268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08098__A2 (.I(_02416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08098__B (.I(_02417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08099__A2 (.I(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08101__A1 (.I(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08101__A2 (.I(_02416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08101__B (.I(_02417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08102__A2 (.I(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08103__A1 (.I(\as2650.stack[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08104__A1 (.I(_02276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08104__A2 (.I(_02416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08104__B (.I(_02417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08105__A2 (.I(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08106__I (.I(_02412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08107__I (.I(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08108__A1 (.I(\as2650.stack[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08109__A1 (.I(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08109__A2 (.I(_02416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08109__B (.I(_02417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08110__A1 (.I(_01884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08111__A1 (.I(\as2650.stack[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08112__I (.I(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08113__A2 (.I(_02428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08114__A1 (.I(_01896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08116__A2 (.I(_02428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08117__A1 (.I(_01909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08119__A2 (.I(_02428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08120__A1 (.I(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08122__A2 (.I(_02428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08123__I (.I(_02412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08124__A1 (.I(_02377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08125__I (.I(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08127__A1 (.I(_02381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08129__A1 (.I(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08131__A1 (.I(_02386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08133__A1 (.I(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08135__A1 (.I(_02390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08137__A1 (.I(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08139__A1 (.I(_02007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08139__A2 (.I(_02253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08141__I (.I(_02446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08143__I (.I(_02446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08144__A2 (.I(_02449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08145__I (.I(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08146__A1 (.I(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08146__A2 (.I(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08147__I (.I(_02452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08148__A2 (.I(_02299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08150__I (.I(_02455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08151__A1 (.I(_02377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08152__I (.I(_02446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08154__A1 (.I(_02381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08156__A1 (.I(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08158__A1 (.I(_02386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08161__I (.I(_02455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08162__A1 (.I(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08163__A1 (.I(\as2650.stack[8][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08164__A1 (.I(_02390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08166__A1 (.I(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08167__I (.I(_02452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08168__A2 (.I(_02299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08169__I (.I(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08171__I (.I(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08172__A2 (.I(_02470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08173__A2 (.I(_02318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08175__I (.I(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08176__A1 (.I(_02377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08177__I (.I(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08179__A1 (.I(_02381_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08181__A1 (.I(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08183__A1 (.I(_02386_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08186__I (.I(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08187__A1 (.I(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08189__A1 (.I(_02390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08191__A1 (.I(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08192__I (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08193__I (.I(_02484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08195__A2 (.I(_01928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08195__A3 (.I(_00981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08195__A4 (.I(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08196__A1 (.I(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08197__A2 (.I(_00975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08197__A4 (.I(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08199__A1 (.I(_00832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08200__A1 (.I(_02490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08201__A1 (.I(_00533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08201__A3 (.I(_00571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08203__A2 (.I(_00482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08206__A3 (.I(_02497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08207__A3 (.I(_02498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08208__A1 (.I(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08209__A1 (.I(_00995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08210__A2 (.I(_00502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08211__A1 (.I(_00529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08214__A2 (.I(_00576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08217__A2 (.I(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08218__A1 (.I(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08218__A2 (.I(_02506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08219__A1 (.I(_02504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08220__A1 (.I(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08221__I (.I(_00571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08222__A2 (.I(_00673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08224__I (.I(_02515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08225__A3 (.I(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08226__A2 (.I(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08228__A2 (.I(_00954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08228__B1 (.I(_02519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08229__A1 (.I(_00749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08230__A1 (.I(_00832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08231__A1 (.I(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08231__A3 (.I(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08232__I (.I(_02523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08234__A1 (.I(_01061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08234__A3 (.I(_00981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08234__A4 (.I(_02525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08235__A1 (.I(_02520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08235__A2 (.I(_02521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08237__A1 (.I(_00749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08237__A2 (.I(_00561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08238__A1 (.I(_00936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08240__A1 (.I(_00836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08240__A3 (.I(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08241__A2 (.I(_00965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08241__A3 (.I(_02525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08245__I (.I(_02536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08246__A2 (.I(_00681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08247__A1 (.I(_00523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08247__A2 (.I(_02537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08247__B (.I(_02538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08248__A2 (.I(_00533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08248__A3 (.I(_00981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08248__A4 (.I(_01787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08249__A2 (.I(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08249__A3 (.I(_02525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08250__A1 (.I(_01108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08251__A1 (.I(_00726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08252__A1 (.I(_02537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08256__I (.I(_02547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08257__I (.I(_00535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08258__A1 (.I(_02146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08258__A2 (.I(_02549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08259__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08260__I (.I(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08262__I (.I(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08263__I (.I(_02554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08264__A1 (.I(_05725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08264__A2 (.I(_02339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08266__A1 (.I(_02554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08266__A2 (.I(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08268__I (.I(_02559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08269__I (.I(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08270__I (.I(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08271__A1 (.I(_02484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08271__A2 (.I(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08271__C (.I(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08274__I (.I(_02565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08275__I (.I(_02566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08276__A1 (.I(_02550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08276__B (.I(_02567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08277__A1 (.I(_02548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08279__C (.I(_02570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08280__I (.I(_02186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08282__I (.I(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08284__I (.I(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08285__A1 (.I(\as2650.stack[6][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08285__A2 (.I(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08286__A2 (.I(_02191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08288__I (.I(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08289__A1 (.I(_02571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08290__I (.I(_02198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08291__I (.I(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08293__A1 (.I(_02580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08294__I (.I(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08296__A1 (.I(_02583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08297__I (.I(_02211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08299__A1 (.I(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08300__I (.I(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08303__I (.I(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08304__A1 (.I(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08305__I (.I(_02225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08307__A1 (.I(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08308__I (.I(_02232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08310__A1 (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08312__I (.I(_02595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08314__I (.I(_02595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08315__A1 (.I(\as2650.stack[5][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08316__A2 (.I(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08318__I (.I(_02601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08319__A1 (.I(_02571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08320__I (.I(_02595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08322__A1 (.I(_02580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08324__A1 (.I(_02583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08326__A1 (.I(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08329__I (.I(_02601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08330__A1 (.I(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08331__A1 (.I(\as2650.stack[5][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08332__A1 (.I(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08333__A1 (.I(\as2650.stack[5][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08334__A1 (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08336__I (.I(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08338__I (.I(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08339__A1 (.I(\as2650.stack[4][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08341__A2 (.I(_02617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08343__I (.I(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08344__A1 (.I(_02571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08345__I (.I(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08347__A1 (.I(_02580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08349__A1 (.I(_02583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08351__A1 (.I(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08354__I (.I(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08355__A1 (.I(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08357__A1 (.I(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08359__A1 (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08360__I (.I(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08363__A2 (.I(_01785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08363__A3 (.I(_02399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08364__I (.I(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08366__A1 (.I(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08367__A1 (.I(_02630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08367__A2 (.I(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08367__B2 (.I(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08368__I (.I(_01846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08369__A1 (.I(\as2650.stack[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08370__I (.I(_02293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08371__I (.I(_02301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08372__A1 (.I(_02268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08372__A2 (.I(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08372__B (.I(_02640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08373__A1 (.I(_02637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08373__A2 (.I(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08374__I (.I(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08376__A1 (.I(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08376__A2 (.I(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08376__B (.I(_02640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08377__A1 (.I(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08377__A2 (.I(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08378__I (.I(_01873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08380__A1 (.I(_02276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08380__A2 (.I(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08380__B (.I(_02640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08381__A1 (.I(_02645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08381__A2 (.I(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08382__I (.I(_01883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08383__I (.I(_02301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08384__I (.I(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08385__A1 (.I(\as2650.stack[12][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08386__A1 (.I(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08386__A2 (.I(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08386__B (.I(_02640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08387__A1 (.I(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08388__I (.I(_01895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08390__A2 (.I(_02296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08391__A1 (.I(_02653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08392__I (.I(_01908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08393__A1 (.I(\as2650.stack[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08394__A2 (.I(_02296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08395__A1 (.I(_02656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08396__I (.I(_01918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08398__A2 (.I(_02296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08399__A1 (.I(_02659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08400__A2 (.I(_02617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08401__I (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08403__I (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08404__A1 (.I(\as2650.stack[3][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08404__A2 (.I(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08405__I (.I(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08406__A2 (.I(_02318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08408__I (.I(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08409__A1 (.I(_02571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08410__I (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08412__A1 (.I(_02580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08414__A1 (.I(_02583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08416__A1 (.I(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08419__I (.I(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08420__A1 (.I(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08422__A1 (.I(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08424__A1 (.I(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08425__I (.I(_02186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08427__I (.I(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08429__I (.I(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08430__A1 (.I(\as2650.stack[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08430__A2 (.I(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08431__A2 (.I(_02191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08431__A3 (.I(_02407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08433__I (.I(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08434__A1 (.I(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08435__I (.I(_02198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08436__I (.I(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08438__A1 (.I(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08439__I (.I(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08441__A1 (.I(_02692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08442__I (.I(_02211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08443__A1 (.I(\as2650.stack[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08444__A1 (.I(_02694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08445__I (.I(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08448__I (.I(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08449__A1 (.I(_02696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08450__I (.I(_02225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08451__A1 (.I(\as2650.stack[2][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08452__A1 (.I(_02700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08453__I (.I(_02232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08455__A1 (.I(_02702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08457__I (.I(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08459__I (.I(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08460__A1 (.I(\as2650.stack[1][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08460__A2 (.I(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08461__A2 (.I(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08461__A3 (.I(_02407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08463__I (.I(_02710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08464__A1 (.I(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08465__I (.I(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08467__A1 (.I(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08469__A1 (.I(_02692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08470__A1 (.I(\as2650.stack[1][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08471__A1 (.I(_02694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08474__I (.I(_02710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08475__A1 (.I(_02696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08477__A1 (.I(_02700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08479__A1 (.I(_02702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08480__A2 (.I(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08481__I (.I(_02721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08483__I (.I(_02721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08484__A2 (.I(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08485__A2 (.I(_01778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08485__A3 (.I(_02318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08487__I (.I(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08488__A1 (.I(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08489__I (.I(_02721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08491__A1 (.I(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08493__A1 (.I(_02692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08495__A1 (.I(_02694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08498__I (.I(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08499__A1 (.I(_02696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08500__A1 (.I(\as2650.stack[15][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08501__A1 (.I(_02700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08503__A1 (.I(_02702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08506__A1 (.I(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08506__A2 (.I(_02739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08508__B1 (.I(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08511__A1 (.I(_00944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08511__B2 (.I(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08512__A1 (.I(_00782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08512__A2 (.I(_00894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08512__A3 (.I(_00967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08512__A4 (.I(_00544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08515__I (.I(_00982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08516__I (.I(_02739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08517__A2 (.I(_00571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08517__A3 (.I(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08517__B1 (.I(_02749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08517__B2 (.I(_02750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08518__A1 (.I(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08519__A2 (.I(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08520__A1 (.I(_00913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08520__A3 (.I(_02749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08520__A4 (.I(_01787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08521__A1 (.I(_00625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08521__B (.I(_00904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08523__A1 (.I(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08523__A2 (.I(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08524__A2 (.I(_00813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08524__B (.I(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08525__A1 (.I(_00502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08525__C (.I(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08527__I (.I(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08529__A3 (.I(_00671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08530__B1 (.I(_02761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08530__B2 (.I(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08532__A1 (.I(_00791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08532__A3 (.I(_01063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08532__B1 (.I(_02761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08535__A1 (.I(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08535__A3 (.I(_00822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08536__A1 (.I(_00913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08536__A2 (.I(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08536__A3 (.I(_02761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08536__A4 (.I(_02339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08537__A1 (.I(_00804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08537__A3 (.I(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08538__A1 (.I(_00815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08540__A4 (.I(_00700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08541__A1 (.I(_01108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08541__A2 (.I(_00826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08541__A3 (.I(_02498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08542__A2 (.I(_00813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08545__A1 (.I(_01271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08545__A2 (.I(_01208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08545__A3 (.I(_01053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08546__A1 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08546__A2 (.I(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08546__A3 (.I(_01420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08546__A4 (.I(_01324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08548__I (.I(_01703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08549__A1 (.I(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08549__A2 (.I(_00817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08550__I (.I(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08551__A1 (.I(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08551__A2 (.I(_00956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08551__A3 (.I(_01697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08553__A1 (.I(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08553__A2 (.I(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08553__A3 (.I(_01304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08553__A4 (.I(_01373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08554__A1 (.I(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08555__A1 (.I(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08555__A2 (.I(_01694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08556__A1 (.I(_01514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08556__A2 (.I(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08562__A1 (.I(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08564__A1 (.I(_01350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08564__A2 (.I(_01180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08564__A3 (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08576__A1 (.I(_01845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08577__A1 (.I(_02798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08578__A1 (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08580__A1 (.I(_00795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08581__A1 (.I(_00538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08582__I (.I(_00839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08583__I (.I(_01942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08584__I (.I(_02817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08587__I (.I(_01953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08588__A1 (.I(\as2650.stack[8][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08588__B2 (.I(\as2650.stack[9][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08591__A1 (.I(\as2650.stack[11][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08591__A2 (.I(_02824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08591__B1 (.I(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08591__B2 (.I(\as2650.stack[10][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08596__A1 (.I(\as2650.stack[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08596__B2 (.I(\as2650.stack[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08597__A1 (.I(\as2650.stack[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08597__B2 (.I(\as2650.stack[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08598__A1 (.I(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08602__A2 (.I(_02835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08602__B1 (.I(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08605__A1 (.I(\as2650.stack[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08605__A2 (.I(_02837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08605__B1 (.I(_02838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08606__A1 (.I(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08607__A1 (.I(\as2650.stack[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08607__A2 (.I(_02837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08607__B1 (.I(_02838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08608__I (.I(_01953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08609__A2 (.I(_02835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08609__B2 (.I(\as2650.stack[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08610__A1 (.I(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08611__B (.I(_01943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08613__I (.I(_02846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08614__I (.I(_00897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08615__I (.I(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08616__I (.I(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08617__I (.I(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08618__I (.I(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08619__I (.I(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08620__I (.I(_02853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08621__A1 (.I(_02850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08621__A2 (.I(_02554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08621__A3 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08622__I (.I(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08623__I (.I(_02856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08624__I (.I(_01216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08625__I (.I(_01265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08626__I (.I(_02859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08627__I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08628__I (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08629__I (.I(_02862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08630__I (.I(_02863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08631__I (.I(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08632__A1 (.I(_02857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08632__A2 (.I(_02858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08632__A3 (.I(_02860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08632__A4 (.I(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08633__B (.I(_00851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08637__A1 (.I(_01921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08637__B (.I(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08638__A1 (.I(_01911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08638__A2 (.I(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08639__A1 (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08639__A2 (.I(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08639__C (.I(_02750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08640__A1 (.I(_02853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08641__A2 (.I(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08642__I (.I(_01061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08643__I (.I(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08644__A1 (.I(_00536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08646__A1 (.I(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08646__A2 (.I(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08648__A1 (.I(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08650__I (.I(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08651__I (.I(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08652__A1 (.I(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08652__A2 (.I(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08652__A3 (.I(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08653__A1 (.I(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08653__A2 (.I(_05851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08654__I (.I(_00897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08655__A1 (.I(_00963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08657__I (.I(_02490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08658__A1 (.I(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08659__A1 (.I(_00807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08660__A2 (.I(_02778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08660__B (.I(_00883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08661__A1 (.I(_02778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08662__A2 (.I(_02778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08662__B (.I(_00846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08663__I (.I(_01067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08664__A1 (.I(_02896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08664__A2 (.I(_00817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08664__C (.I(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08665__A1 (.I(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08667__B (.I(_00553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08668__I (.I(_00529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08670__I (.I(_02902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08672__I (.I(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08673__A1 (.I(_00849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08673__A2 (.I(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08674__A1 (.I(_02862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08674__A2 (.I(_01261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08674__B1 (.I(_01072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08674__B2 (.I(_01214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08676__A1 (.I(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08676__A2 (.I(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08676__B1 (.I(_01211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08676__B2 (.I(_01265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08678__A1 (.I(_00943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08679__A1 (.I(_02910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08679__A2 (.I(_01067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08679__B1 (.I(_01522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08679__B2 (.I(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08679__C (.I(_02911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08680__A1 (.I(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08680__A2 (.I(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08680__B1 (.I(_01224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08680__B2 (.I(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08682__I (.I(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08683__A2 (.I(_01215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08683__B1 (.I(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08683__B2 (.I(_05735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08684__A1 (.I(_01007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08684__A2 (.I(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08684__B1 (.I(_01536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08684__B2 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08685__A1 (.I(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08685__A2 (.I(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08685__B1 (.I(_02862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08685__B2 (.I(_01872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08686__A1 (.I(_05727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08686__A2 (.I(_02910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08686__B1 (.I(_01265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08686__B2 (.I(_01861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08687__A1 (.I(_02911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08688__A1 (.I(_01350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08688__A2 (.I(_00625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08688__A3 (.I(_00469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08690__I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08691__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08693__A2 (.I(_02925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08693__B1 (.I(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08693__B2 (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08694__A1 (.I(_02173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08694__A2 (.I(_01079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08694__B1 (.I(_01215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08694__B2 (.I(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08695__A2 (.I(_01328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08695__B1 (.I(_01536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08695__B2 (.I(_02484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08696__A1 (.I(_02923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08696__A2 (.I(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08696__B2 (.I(_00848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08697__A1 (.I(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08698__A1 (.I(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08699__I (.I(_02910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08700__A2 (.I(_02932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08701__A1 (.I(_02497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08703__A1 (.I(_00793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08703__B (.I(_02345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08705__I (.I(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08708__I (.I(_00602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08710__A1 (.I(_02942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08710__A2 (.I(_02902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08711__A1 (.I(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08712__A2 (.I(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08713__I (.I(_01942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08714__A2 (.I(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08714__B2 (.I(\as2650.stack[9][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08715__A1 (.I(\as2650.stack[11][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08715__A2 (.I(_02837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08715__B1 (.I(_02838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08716__A1 (.I(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08719__A1 (.I(\as2650.stack[15][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08719__A2 (.I(_02951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08719__B1 (.I(_02838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08720__A2 (.I(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08721__A1 (.I(_02950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08723__A2 (.I(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08725__A1 (.I(\as2650.stack[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08725__A2 (.I(_02951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08725__B1 (.I(_02957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08725__B2 (.I(\as2650.stack[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08726__A1 (.I(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08727__A1 (.I(\as2650.stack[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08727__A2 (.I(_02951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08727__B1 (.I(_02957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08727__B2 (.I(\as2650.stack[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08729__I (.I(_01953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08730__A1 (.I(\as2650.stack[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08730__A2 (.I(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08730__B1 (.I(_02962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08730__B2 (.I(\as2650.stack[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08731__A1 (.I(_02950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08732__B (.I(_02817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08733__A1 (.I(_02946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08734__A1 (.I(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08734__A2 (.I(_02966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08735__A1 (.I(_02778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08739__A2 (.I(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08741__A1 (.I(\as2650.stack[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08742__I (.I(_01839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08743__A1 (.I(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08744__A1 (.I(_02630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08744__B2 (.I(_02975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08745__A1 (.I(\as2650.stack[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08746__I (.I(_01857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08747__I (.I(_02721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08748__I (.I(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08749__A1 (.I(_02977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08750__A1 (.I(_02637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08751__A1 (.I(\as2650.stack[15][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08752__I (.I(_01869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08753__A1 (.I(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08754__A1 (.I(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08755__A1 (.I(\as2650.stack[15][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08756__I (.I(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08757__A1 (.I(_02985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08758__A1 (.I(_02645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08759__I (.I(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08761__A1 (.I(\as2650.stack[15][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08762__I (.I(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08763__A1 (.I(_02990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08764__A1 (.I(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08765__A1 (.I(\as2650.stack[15][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08766__I (.I(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08767__A1 (.I(_02993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08767__A2 (.I(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08768__A1 (.I(_02653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08769__A1 (.I(\as2650.stack[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08770__I (.I(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08771__A1 (.I(_02996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08771__A2 (.I(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08772__A1 (.I(_02656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08773__A1 (.I(\as2650.stack[15][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08774__I (.I(_01924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08775__A1 (.I(_02999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08775__A2 (.I(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08776__A1 (.I(_02659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08779__A1 (.I(_02250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08780__I (.I(_03003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08781__A1 (.I(\as2650.stack[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08782__A1 (.I(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08783__A1 (.I(_02630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08783__B2 (.I(_03006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08784__A1 (.I(\as2650.stack[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08785__I (.I(_02446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08786__I (.I(_02455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08787__A1 (.I(_02977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08788__A1 (.I(_02637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08789__A1 (.I(\as2650.stack[8][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08790__A1 (.I(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08791__A1 (.I(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08792__A1 (.I(\as2650.stack[8][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08793__A1 (.I(_02985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08794__A1 (.I(_02645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08795__I (.I(_02455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08796__I (.I(_03003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08797__A1 (.I(\as2650.stack[8][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08798__A1 (.I(_02990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08799__A1 (.I(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08800__A1 (.I(\as2650.stack[8][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08801__A1 (.I(_02993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08801__A2 (.I(_02449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08802__A1 (.I(_02653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08803__A1 (.I(\as2650.stack[8][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08804__A1 (.I(_02996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08804__A2 (.I(_02449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08805__A1 (.I(_02656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08807__A1 (.I(_02999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08807__A2 (.I(_02449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08808__A1 (.I(_02659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08812__A1 (.I(_02250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08812__A2 (.I(_02253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08812__A3 (.I(_03027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08813__I (.I(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08814__A1 (.I(\as2650.stack[11][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08815__A1 (.I(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08816__A1 (.I(_02630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08817__A1 (.I(\as2650.stack[11][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08818__I (.I(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08819__I (.I(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08820__A1 (.I(_02977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08821__A1 (.I(_02637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08822__A1 (.I(\as2650.stack[11][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08823__A1 (.I(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08824__A1 (.I(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08825__A1 (.I(\as2650.stack[11][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08826__A1 (.I(_02985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08827__A1 (.I(_02645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08828__I (.I(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08829__I (.I(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08830__A1 (.I(\as2650.stack[11][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08831__A1 (.I(_02990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08832__A1 (.I(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08833__A1 (.I(\as2650.stack[11][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08834__A1 (.I(_02993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08834__A2 (.I(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08835__A1 (.I(_02653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08836__A1 (.I(\as2650.stack[11][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08837__A1 (.I(_02996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08837__A2 (.I(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08838__A1 (.I(_02656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08839__A1 (.I(\as2650.stack[11][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08840__A1 (.I(_02999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08840__A2 (.I(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08841__A1 (.I(_02659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08842__I (.I(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08846__I (.I(_03053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08847__A1 (.I(\as2650.stack[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08848__A1 (.I(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08849__A1 (.I(_03050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08849__A2 (.I(_03052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08849__B2 (.I(_03056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08850__I (.I(_01846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08852__I (.I(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08853__I (.I(_02710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08854__A1 (.I(_02977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08854__A2 (.I(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08854__B (.I(_03060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08855__A1 (.I(_03057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08855__A2 (.I(_03052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08856__I (.I(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08858__A1 (.I(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08858__A2 (.I(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08858__B (.I(_03060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08859__A1 (.I(_03062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08859__A2 (.I(_03052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08860__I (.I(_01873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08862__A1 (.I(_02985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08862__A2 (.I(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08862__B (.I(_03060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08863__A1 (.I(_03065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08863__A2 (.I(_03052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08864__I (.I(_01883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08865__I (.I(_02710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08866__I (.I(_03053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08868__A1 (.I(_02990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08868__A2 (.I(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08868__B (.I(_03060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08869__A1 (.I(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08870__I (.I(_01895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08872__A1 (.I(_02993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08872__A2 (.I(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08873__A1 (.I(_03073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08874__I (.I(_01908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08876__A1 (.I(_02996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08876__A2 (.I(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08877__A1 (.I(_03076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08878__I (.I(_01918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08880__A1 (.I(_02999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08880__A2 (.I(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08881__A1 (.I(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08882__A1 (.I(_05781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08884__A1 (.I(_00814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08884__A2 (.I(_01022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08884__A3 (.I(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08885__I (.I(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08886__A1 (.I(_01007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08886__A2 (.I(_00475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08887__A2 (.I(_03086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08890__A4 (.I(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08891__A1 (.I(_00622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08891__A2 (.I(_01014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08891__A3 (.I(_01017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08892__A1 (.I(_01007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08892__A2 (.I(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08893__I (.I(_03092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08894__A1 (.I(_01028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08894__A2 (.I(_01029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08894__A3 (.I(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08896__A1 (.I(_00673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08896__A3 (.I(_01004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08897__I (.I(_03096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08900__A3 (.I(_03090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08901__I (.I(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08902__A1 (.I(_00989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08903__I (.I(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08905__I (.I(_03090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08906__I (.I(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08907__A1 (.I(_00671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08907__A3 (.I(_03086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08909__I (.I(_01079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08911__I (.I(_03096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08912__A1 (.I(_00455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08913__A1 (.I(_03109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08914__A3 (.I(_03086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08916__A1 (.I(_01072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08917__I (.I(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08920__A1 (.I(_01054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08921__I (.I(_03090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08923__A1 (.I(_01094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08925__A1 (.I(_01051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08926__I (.I(_03092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08928__I0 (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08929__A1 (.I(_01008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08929__A2 (.I(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08930__A1 (.I(_00978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08931__A1 (.I(_00989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08931__A2 (.I(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08931__C (.I(_00599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08932__I (.I(_03131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08935__I (.I(_03134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08936__A1 (.I(_01142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08936__A2 (.I(_01146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08937__A2 (.I(_03128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08938__I (.I(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08940__A1 (.I(_01032_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08940__A3 (.I(_03086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08941__I (.I(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08943__A1 (.I(_00454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08944__A1 (.I(_01216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08946__A1 (.I(_01212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08947__A1 (.I(_00953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08947__A2 (.I(_01061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08949__A1 (.I(_01224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08950__A1 (.I(_01209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08951__A1 (.I(_01206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08953__A1 (.I(_01199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08954__I0 (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08956__A2 (.I(_03153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08957__I (.I(_01072_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08958__A1 (.I(_00657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08958__A2 (.I(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08958__A3 (.I(_01004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08958__A4 (.I(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08959__I (.I(_03156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08960__A1 (.I(_00953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08961__A1 (.I(_00450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08961__A2 (.I(_03156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08962__A1 (.I(_02859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08963__A1 (.I(_00434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08964__A1 (.I(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08965__I0 (.I(_01272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08967__A1 (.I(_01260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08968__A1 (.I(_01254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08969__A1 (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08972__A2 (.I(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08973__A1 (.I(_00452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08974__A1 (.I(_02863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08975__A1 (.I(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08977__A1 (.I(_01212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08978__A1 (.I(_01325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08979__A1 (.I(_01323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08982__A1 (.I(_01343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08983__I0 (.I(_01373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08984__A1 (.I(_01230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08984__A2 (.I(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08985__A1 (.I(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08985__A2 (.I(_03181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08987__A2 (.I(_03180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08988__I (.I(_03181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08989__I (.I(_03131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08990__A1 (.I(\as2650.r123_2[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08991__A1 (.I(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08993__I (.I(_03090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08994__A1 (.I(_00437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08995__A1 (.I(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08996__A1 (.I(_00425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08997__A1 (.I(_01262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__08998__A1 (.I(_01420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09000__A1 (.I(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09001__A1 (.I(_01413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09003__A1 (.I(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09005__A2 (.I(_03200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09008__I (.I(_01535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09009__A1 (.I(_03203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09010__A1 (.I(_00428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09011__A1 (.I(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09012__A1 (.I(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09013__A1 (.I(_02146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09014__A1 (.I(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09016__A1 (.I(_01526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09018__A1 (.I(_01514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09019__A1 (.I(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09019__B2 (.I(\as2650.r123_2[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09020__A2 (.I(_03213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09021__A1 (.I(_00424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09022__A1 (.I(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09023__A1 (.I(_02896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09024__A1 (.I(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09025__A1 (.I(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09026__A1 (.I(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09028__A1 (.I(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09030__A1 (.I(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09031__A1 (.I(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09031__A2 (.I(_03134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09031__B2 (.I(\as2650.r123_2[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09032__A2 (.I(_03224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09033__A1 (.I(\as2650.r123_2[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09034__A1 (.I(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09035__I (.I(_01694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09036__I0 (.I(_00421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09036__I1 (.I(_00602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09039__A1 (.I(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09040__A1 (.I(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09041__A1 (.I(_01713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09043__A1 (.I(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09045__A1 (.I(_03228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09046__A2 (.I(_03238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09049__A2 (.I(_00984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09050__A1 (.I(_03134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09052__A1 (.I(_01230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09052__A2 (.I(_00942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09054__A1 (.I(_01990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09057__A1 (.I(_01142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09058__A1 (.I(_05763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09060__B2 (.I(_03128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09061__A1 (.I(_05718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09064__I0 (.I(\as2650.r123_2[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09064__I1 (.I(_03252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09064__S (.I(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09066__A1 (.I(_02042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09067__A1 (.I(_01850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09068__B2 (.I(_03153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09069__I1 (.I(_03259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09069__S (.I(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09071__A1 (.I(_02065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09072__A1 (.I(_01865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09073__B2 (.I(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09074__I1 (.I(_03263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09074__S (.I(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09078__A1 (.I(_02095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09079__A1 (.I(_02097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09081__B2 (.I(_03180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09082__I0 (.I(\as2650.r123_2[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09082__I1 (.I(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09082__S (.I(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09084__A1 (.I(_02118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09085__A1 (.I(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09086__B2 (.I(_03200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09088__I1 (.I(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09090__A1 (.I(_02144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09091__A1 (.I(_02146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09092__B2 (.I(_03213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09095__A1 (.I(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09096__A1 (.I(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09097__B2 (.I(_03224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09098__I0 (.I(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09100__I (.I(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09101__A1 (.I(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09102__A1 (.I(_03238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09106__I (.I(_03289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09107__A1 (.I(_02406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09108__A1 (.I(_02250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09108__A2 (.I(_03027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09111__I (.I(_01839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09112__A1 (.I(_03295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09113__A1 (.I(_03050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09113__B2 (.I(_03296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09114__A1 (.I(\as2650.stack[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09115__I (.I(_01857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09116__I (.I(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09117__I (.I(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09118__A2 (.I(_03299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09118__B (.I(_03300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09119__A1 (.I(_03057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09120__A1 (.I(\as2650.stack[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09121__I (.I(_01869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09122__A2 (.I(_03299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09122__B (.I(_03300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09123__A1 (.I(_03062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09125__I (.I(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09126__A2 (.I(_03299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09126__B (.I(_03300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09127__A1 (.I(_03065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09128__I (.I(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09130__A2 (.I(_03309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09131__I (.I(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09132__A2 (.I(_03299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09132__B (.I(_03300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09133__A1 (.I(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09133__A2 (.I(_03308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09134__A1 (.I(\as2650.stack[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09134__A2 (.I(_03309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09135__I (.I(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09136__A2 (.I(_02470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09136__B (.I(_03289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09137__A1 (.I(_03073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09137__A2 (.I(_03308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09138__A1 (.I(\as2650.stack[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09138__A2 (.I(_03309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09139__I (.I(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09140__A2 (.I(_02470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09140__B (.I(_03289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09141__A1 (.I(_03076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09141__A2 (.I(_03308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09142__A1 (.I(\as2650.stack[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09142__A2 (.I(_03309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09143__I (.I(_01924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09144__A2 (.I(_02470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09144__B (.I(_03289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09145__A1 (.I(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09145__A2 (.I(_03308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09164__A1 (.I(_05786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09164__A3 (.I(_05765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09165__B2 (.I(_05786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09167__A1 (.I(_05854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09175__A1 (.I(_05808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09175__A2 (.I(_01733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09177__A1 (.I(_05797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09178__A2 (.I(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09184__A1 (.I(_00947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09186__A1 (.I(_00947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09186__B (.I(_03134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09186__C (.I(_00909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09189__A1 (.I(_03322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09189__A2 (.I(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09189__B1 (.I(_03361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09189__B2 (.I(_03128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09197__A2 (.I(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09204__A1 (.I(_05808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09207__A1 (.I(\as2650.r0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09207__A3 (.I(_05765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09208__B2 (.I(\as2650.r0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09210__A1 (.I(\as2650.r0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09215__A2 (.I(_01733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09216__A1 (.I(_05787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09216__A2 (.I(_01640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09225__A1 (.I(_03153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09225__B1 (.I(_03397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09230__A1 (.I(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09230__A2 (.I(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09231__A1 (.I(_01420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09231__A2 (.I(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09236__A1 (.I(_05855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09236__A2 (.I(_01640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09241__A1 (.I(_05809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09243__A1 (.I(_05807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09244__A1 (.I(_05758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09248__A1 (.I(_05797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09257__A1 (.I(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09257__B1 (.I(_03429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09264__A1 (.I(_05758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09264__A2 (.I(_01724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09271__A1 (.I(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09273__A2 (.I(_05767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09276__A1 (.I(_05787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09287__A1 (.I(_03180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09287__B1 (.I(_03458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09297__A1 (.I(_05855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09298__A2 (.I(_05767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09304__A1 (.I(_03464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09305__A1 (.I(_03461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09308__A1 (.I(_03200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09308__B1 (.I(_03477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09309__A1 (.I(_03464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09310__A1 (.I(_03461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09315__I (.I(_05767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09316__A1 (.I(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09316__A2 (.I(_03486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09316__B1 (.I(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09317__A3 (.I(_03486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09317__A4 (.I(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09319__A1 (.I(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09326__A1 (.I(_03213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09326__A2 (.I(_03361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09326__B1 (.I(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09326__B2 (.I(_03322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09327__A1 (.I(_01703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09330__A1 (.I(_03486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09331__S (.I(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09334__A1 (.I(_03224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09334__A2 (.I(_03361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09334__B1 (.I(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09334__B2 (.I(_03322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09339__A1 (.I(_03238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09339__A2 (.I(_03361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09339__B1 (.I(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09339__B2 (.I(_03322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09341__I (.I(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09343__A2 (.I(_03027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09345__A1 (.I(\as2650.stack[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09346__A1 (.I(_03295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09347__A1 (.I(_03050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09347__B2 (.I(_03514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09348__A1 (.I(\as2650.stack[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09349__I (.I(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09350__I (.I(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09351__A2 (.I(_03516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09351__B (.I(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09352__A1 (.I(_03057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09353__A1 (.I(\as2650.stack[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09354__A2 (.I(_03516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09354__B (.I(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09355__A1 (.I(_03062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09357__A2 (.I(_03516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09357__B (.I(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09358__A1 (.I(_03065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09359__I (.I(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09361__A1 (.I(\as2650.stack[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09362__A2 (.I(_03516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09362__B (.I(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09363__A1 (.I(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09363__A2 (.I(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09364__A1 (.I(\as2650.stack[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09365__A2 (.I(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09365__B (.I(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09366__A1 (.I(_03073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09366__A2 (.I(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09367__A1 (.I(\as2650.stack[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09368__A2 (.I(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09368__B (.I(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09369__A1 (.I(_03076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09369__A2 (.I(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09370__A1 (.I(\as2650.stack[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09371__A2 (.I(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09371__B (.I(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09372__A1 (.I(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09372__A2 (.I(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09374__I (.I(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09377__A1 (.I(\as2650.stack[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09378__A1 (.I(_03295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09379__A1 (.I(_03050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09379__B2 (.I(_03538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09380__A1 (.I(\as2650.stack[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09381__I (.I(_02595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09382__I (.I(_02601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09383__A2 (.I(_03540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09383__B (.I(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09384__A1 (.I(_03057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09385__A1 (.I(\as2650.stack[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09386__A2 (.I(_03540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09386__B (.I(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09387__A1 (.I(_03062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09388__A1 (.I(\as2650.stack[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09389__A2 (.I(_03540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09389__B (.I(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09390__A1 (.I(_03065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09391__I (.I(_02601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09393__A1 (.I(\as2650.stack[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09394__A2 (.I(_03540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09394__B (.I(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09395__A1 (.I(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09396__A1 (.I(\as2650.stack[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09397__B (.I(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09398__A1 (.I(_03073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09399__A1 (.I(\as2650.stack[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09400__B (.I(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09401__A1 (.I(_03076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09402__A1 (.I(\as2650.stack[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09403__B (.I(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09404__A1 (.I(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09405__I (.I(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09407__I (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09408__A1 (.I(_02399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09411__A1 (.I(_03295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09412__A1 (.I(_03557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09412__B2 (.I(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09413__I (.I(_01845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09415__I (.I(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09416__I (.I(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09417__A2 (.I(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09417__B (.I(_03567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09418__A1 (.I(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09419__I (.I(_01861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09420__A1 (.I(\as2650.stack[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09421__A2 (.I(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09421__B (.I(_03567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09422__A1 (.I(_03569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09423__I (.I(_01872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09425__A2 (.I(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09425__B (.I(_03567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09426__A1 (.I(_03572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09427__I (.I(_01883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09428__I (.I(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09431__A2 (.I(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09431__B (.I(_03567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09435__B (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09436__A1 (.I(_03580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09437__I (.I(_01908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09439__B (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09441__I (.I(_01918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09442__A1 (.I(\as2650.stack[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09443__B (.I(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09447__A2 (.I(_02255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09449__A2 (.I(_03592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09450__A1 (.I(_01840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09451__A1 (.I(_03557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09451__A2 (.I(_03590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09451__B2 (.I(_03594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09452__A1 (.I(\as2650.stack[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09452__A2 (.I(_03592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09453__I (.I(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09454__I (.I(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09455__A2 (.I(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09455__B (.I(_03597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09456__A1 (.I(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09456__A2 (.I(_03590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09457__A1 (.I(\as2650.stack[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09457__A2 (.I(_03592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09458__A1 (.I(_01870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09458__A2 (.I(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09458__B (.I(_03597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09459__A1 (.I(_03569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09459__A2 (.I(_03590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09460__A1 (.I(\as2650.stack[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09460__A2 (.I(_03592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09461__A1 (.I(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09461__A2 (.I(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09461__B (.I(_03597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09462__A1 (.I(_03572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09462__A2 (.I(_03590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09463__I (.I(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09466__A1 (.I(_01892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09466__A2 (.I(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09466__B (.I(_03597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09469__A2 (.I(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09470__A1 (.I(_03580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09472__A2 (.I(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09474__A1 (.I(\as2650.stack[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09475__A2 (.I(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09477__A1 (.I(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09478__A1 (.I(_00599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09478__A2 (.I(_00956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09478__A3 (.I(_00937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09478__A4 (.I(_03613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09479__I (.I(_03614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09481__I (.I(_03614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09483__A1 (.I(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09484__A1 (.I(\as2650.ivec[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09485__A1 (.I(_01851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09486__I0 (.I(\as2650.ivec[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09486__I1 (.I(_02067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09488__I1 (.I(_02098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09490__I (.I(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09491__I1 (.I(_03622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09494__A1 (.I(_01900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09495__I (.I(_01911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09497__A1 (.I(_03625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09498__I0 (.I(\as2650.ivec[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09498__I1 (.I(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09498__S (.I(_03614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09502__A2 (.I(_02255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09504__A2 (.I(_03631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09505__A1 (.I(_01840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09506__A1 (.I(_03557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09506__A2 (.I(_03629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09506__B2 (.I(_03633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09507__A1 (.I(\as2650.stack[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09507__A2 (.I(_03631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09508__I (.I(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09509__I (.I(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09510__A2 (.I(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09510__B (.I(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09511__A1 (.I(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09511__A2 (.I(_03629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09512__A2 (.I(_03631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09513__A1 (.I(_01870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09513__A2 (.I(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09513__B (.I(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09514__A1 (.I(_03569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09514__A2 (.I(_03629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09515__A1 (.I(\as2650.stack[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09515__A2 (.I(_03631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09516__A1 (.I(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09516__A2 (.I(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09516__B (.I(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09517__A1 (.I(_03572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09517__A2 (.I(_03629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09518__I (.I(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09520__A2 (.I(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09521__A1 (.I(_01892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09521__A2 (.I(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09521__B (.I(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09523__A2 (.I(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09524__A2 (.I(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09525__A1 (.I(_03580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09526__A2 (.I(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09527__A2 (.I(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09529__A1 (.I(\as2650.stack[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09529__A2 (.I(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09530__A2 (.I(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09532__A2 (.I(_00681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09533__A1 (.I(_00875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09535__A1 (.I(_00832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09538__A1 (.I(_00466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09538__A2 (.I(_00907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09538__A4 (.I(_03657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09539__A1 (.I(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09540__A2 (.I(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09540__B (.I(_00894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09541__A2 (.I(_03653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09542__I (.I(_02750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09543__I (.I(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09544__A1 (.I(_00642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09544__A2 (.I(_00580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09545__A1 (.I(_00928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09546__I (.I(_03653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09547__A1 (.I(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09547__B (.I(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09549__A1 (.I(_00625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09549__A2 (.I(_00647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09552__A1 (.I(_00804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09553__A1 (.I(_00679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09553__A2 (.I(_00533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09554__A1 (.I(_01033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09554__A2 (.I(_03673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09556__A1 (.I(_00709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09556__A2 (.I(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09556__B (.I(_00837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09557__A1 (.I(_00483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09559__I (.I(_00627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09560__I (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09561__I (.I(_00628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09562__A1 (.I(_03681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09562__A2 (.I(_00844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09563__A1 (.I(_03680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09564__A1 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09564__A2 (.I(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09564__B (.I(_00883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09565__A1 (.I(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09565__A2 (.I(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09566__I (.I(_02525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09567__A1 (.I(_00954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09567__A3 (.I(_03685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09568__A1 (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09568__A2 (.I(_03686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09569__I (.I(_00909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09570__I (.I(_03688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09571__A1 (.I(_01118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09571__A2 (.I(_03686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09571__C (.I(_03689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09572__A1 (.I(_00575_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09572__A2 (.I(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09573__A1 (.I(_00642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09573__A2 (.I(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09576__A1 (.I(_00502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09576__B3 (.I(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09578__A1 (.I(_00967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09578__A2 (.I(_02519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09578__C (.I(_00692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09580__A1 (.I(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09580__A2 (.I(_00675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09580__A3 (.I(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09581__B (.I(_02537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09583__B (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09584__I (.I(_00506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09585__I (.I(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09586__A1 (.I(_00576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09586__A2 (.I(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09587__A1 (.I(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09589__A1 (.I(_00459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09589__A2 (.I(_00715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09589__A4 (.I(_03685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09590__A1 (.I(_00944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09591__A2 (.I(_00822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09591__A3 (.I(_03685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09592__A1 (.I(_02515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09592__A2 (.I(_02519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09593__A1 (.I(_00716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09594__A1 (.I(_02565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09595__A1 (.I(_00946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09596__A1 (.I(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09596__A2 (.I(_00978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09597__A3 (.I(_03685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09599__A2 (.I(_00822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09599__A3 (.I(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09600__A1 (.I(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09600__A2 (.I(_00954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09602__A1 (.I(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09603__A2 (.I(_00654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09607__A2 (.I(_03723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09608__A1 (.I(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09609__A1 (.I(_02523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09611__I (.I(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09613__A2 (.I(_03729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09615__A3 (.I(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09616__A1 (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09616__A2 (.I(_00473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09616__A4 (.I(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09617__A2 (.I(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09618__A2 (.I(_00916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09620__A2 (.I(_00495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09621__A2 (.I(_03736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09622__A2 (.I(_00967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09622__C (.I(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09623__A1 (.I(_00660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09623__A2 (.I(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09624__A1 (.I(_01791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09625__A1 (.I(_01033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09625__A2 (.I(_00873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09625__A4 (.I(_02519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09626__B (.I(_03741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09629__A1 (.I(_02504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09629__A3 (.I(_03719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09630__I (.I(_03746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09632__A2 (.I(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09633__A1 (.I(_00969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09634__I (.I(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09635__I (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09638__I (.I(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09640__I (.I(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09641__A2 (.I(_03109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09644__A1 (.I(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09644__A2 (.I(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09646__A1 (.I(_00830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09646__A2 (.I(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09646__A3 (.I(_00732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09647__A1 (.I(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09647__A2 (.I(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09647__C (.I(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09648__I (.I(_01834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09649__A1 (.I(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09650__A2 (.I(_03766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09651__I (.I(_03109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09652__A1 (.I(_00629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09652__A2 (.I(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09654__A1 (.I(_00629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09656__I (.I(_00699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09657__A1 (.I(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09657__B (.I(_02515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09658__A1 (.I(_03768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09658__B2 (.I(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09659__B (.I(_00718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09660__A2 (.I(_02549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09661__A1 (.I(_03754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09661__A2 (.I(_03764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09662__A2 (.I(_00834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09662__B (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09663__I (.I(_00597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09665__A1 (.I(_00754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09665__A2 (.I(_00770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09667__A2 (.I(_01094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09668__I (.I(_00769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09669__A1 (.I(_02856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09670__A1 (.I(_03768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09671__I (.I(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09673__A1 (.I(_01078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09673__A2 (.I(_01050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09674__I (.I(_01103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09676__A2 (.I(_01051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09678__A2 (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09678__B2 (.I(_03768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09681__B1 (.I(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09681__B2 (.I(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09682__A1 (.I(_00598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09682__A2 (.I(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09683__I (.I(_03673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09684__I (.I(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09685__A1 (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09685__C (.I(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09686__A2 (.I(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09687__A1 (.I(_00777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09688__A1 (.I(_01836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09688__A2 (.I(_03751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09689__I (.I(_03746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09691__A1 (.I(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09691__B (.I(_00883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09692__A2 (.I(_03805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09693__I (.I(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09695__A1 (.I(_00526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09695__A2 (.I(_00708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09697__A1 (.I(_00919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09698__A1 (.I(_00829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09698__A2 (.I(_00732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09699__I (.I(_03814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09700__I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09701__I (.I(_00848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09702__I (.I(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09703__A1 (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09703__A2 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09704__A1 (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09704__A2 (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09705__A2 (.I(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09706__A1 (.I(_00850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09706__A2 (.I(_03821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09707__A2 (.I(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09711__I (.I(_00723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09712__A1 (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09713__A1 (.I(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09714__A1 (.I(_02858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09715__B2 (.I(_00734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09716__I (.I(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09718__A1 (.I(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09718__B2 (.I(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09720__I (.I(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09721__I (.I(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09722__A1 (.I(_01834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09722__A2 (.I(_01078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09723__A2 (.I(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09724__I (.I(_00635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09725__I (.I(_01215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09726__I (.I(_01088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09727__A1 (.I(_01078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09727__A2 (.I(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09729__A2 (.I(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09729__A3 (.I(_01203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09733__A1 (.I(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09734__A2 (.I(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09734__A3 (.I(_01196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09735__A1 (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09735__A2 (.I(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09736__A1 (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09736__A2 (.I(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09737__A1 (.I(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09738__A2 (.I(_03849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09740__B (.I(_03855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09742__I (.I(_02559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09743__A1 (.I(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09743__A2 (.I(_03858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09744__A1 (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09744__C (.I(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09745__A1 (.I(_03809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09745__A2 (.I(_03810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09745__B2 (.I(_03837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09745__C (.I(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09746__A1 (.I(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09746__A2 (.I(_03751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09746__B2 (.I(_02548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09747__I (.I(_00845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09749__A2 (.I(_03862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09751__I (.I(_00907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09752__A1 (.I(_03865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09752__A2 (.I(_03866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09753__I (.I(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09754__A1 (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09754__A2 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09755__A1 (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09755__A2 (.I(_01214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09756__A2 (.I(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09756__B (.I(_03870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09757__A1 (.I(_03869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09757__A2 (.I(_03871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09759__I (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09763__A1 (.I(_01216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09763__A2 (.I(_01206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09764__A1 (.I(_01264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09764__A2 (.I(_01260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09767__A1 (.I(_02860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09767__B (.I(_03881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09769__I (.I(_02925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09772__A1 (.I(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09772__B1 (.I(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09772__B2 (.I(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09773__A1 (.I(_03884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09773__A2 (.I(_01254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09773__A3 (.I(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09774__A1 (.I(_03884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09778__B1 (.I(_03891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09779__S (.I(_00610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09781__A1 (.I(_00716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09781__A2 (.I(_00708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09785__A1 (.I(_02859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09786__A2 (.I(_00631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09787__A1 (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09787__C (.I(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09789__I (.I(_00848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09790__I (.I(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09791__A2 (.I(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09791__B (.I(_03870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09792__A1 (.I(_03869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09792__A2 (.I(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09794__A1 (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09794__B (.I(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09795__A1 (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09798__A1 (.I(_01868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09798__A2 (.I(_03895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09798__B2 (.I(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09800__I (.I(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09801__A1 (.I(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09801__B2 (.I(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09803__A1 (.I(_01868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09803__B2 (.I(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09804__A1 (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09805__A2 (.I(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09806__I (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09807__I (.I(_03920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09808__I (.I(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09809__I (.I(_00875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09812__A1 (.I(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09812__A2 (.I(_00794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09813__I (.I(_03858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09814__A2 (.I(_03927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09815__A1 (.I(_03920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09815__A2 (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09817__A1 (.I(_03920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09817__A2 (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09819__A1 (.I(_01866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09819__A2 (.I(_01264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09820__I (.I(_03869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09821__A2 (.I(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09825__A1 (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09825__A2 (.I(_00604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09826__I (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09827__A1 (.I(net99));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09827__A2 (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09829__A1 (.I(_00928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09830__A1 (.I(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09830__B2 (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09830__C (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09832__A1 (.I(_03921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09832__A2 (.I(_03926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09832__B1 (.I(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09834__A2 (.I(_03871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09837__I (.I(_01328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09838__A1 (.I(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09839__A2 (.I(_01259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09840__A3 (.I(_01259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09842__A2 (.I(_01320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09843__A1 (.I(_01262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09845__A1 (.I(_01328_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09845__A2 (.I(_03958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09846__I (.I(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09847__A2 (.I(_01323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09851__A1 (.I(_03951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09851__B (.I(_03964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09851__C (.I(_00636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09852__C (.I(_02925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09853__A1 (.I(_01251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09853__A2 (.I(_01252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09854__C (.I(_02925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09855__A1 (.I(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09856__A1 (.I(_02863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09856__A2 (.I(_01343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09857__A1 (.I(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09859__A2 (.I(_03970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09859__C (.I(_03972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09860__B (.I(_00766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09861__A2 (.I(_00770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09862__B (.I(_00610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09863__A1 (.I(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09865__I (.I(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09866__A1 (.I(_03681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09867__I (.I(_00969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09868__I (.I(_03981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09869__A1 (.I(_03921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09871__A1 (.I(net98));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09873__I (.I(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09874__I (.I(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09875__I (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09876__A1 (.I(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09876__A2 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09880__B (.I(_00597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09883__A2 (.I(_01412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09887__A2 (.I(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09888__A2 (.I(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09889__A1 (.I(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09890__I (.I(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09891__A2 (.I(_01415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09892__A2 (.I(_01323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09894__B (.I(_01088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09896__A1 (.I(_04003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09897__B2 (.I(_00635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09899__B (.I(_04011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09900__B2 (.I(_00598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09901__I (.I(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09902__I (.I(_04014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09903__A1 (.I(_00874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09904__I (.I(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09906__I (.I(_00630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09907__I (.I(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09908__A1 (.I(_00630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09908__A2 (.I(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09909__A2 (.I(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09909__B (.I(_04020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09910__A1 (.I(_00724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09910__C (.I(_00733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09911__I (.I(_02932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09914__A1 (.I(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09914__A2 (.I(_04026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09915__A2 (.I(_00850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09915__B (.I(_03814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09917__A1 (.I(_04015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09917__A2 (.I(_03895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09917__B1 (.I(_04017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09919__A1 (.I(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09919__B2 (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09920__I (.I(_02547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09921__A1 (.I(_01889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09921__B2 (.I(_04033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09923__A1 (.I(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09925__I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09927__A1 (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09927__A2 (.I(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09929__A1 (.I(_04014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09929__A2 (.I(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09931__A1 (.I(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09931__A2 (.I(_04042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09932__A1 (.I(_04037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09932__A2 (.I(_04038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09933__I (.I(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09935__A1 (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09937__I (.I(_04048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09938__A1 (.I(_04045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09938__C2 (.I(_04037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09939__B2 (.I(_00734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09940__A1 (.I(_01903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09940__A2 (.I(_03926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09940__B1 (.I(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09941__A2 (.I(_01413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09942__A2 (.I(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09943__A1 (.I(_03203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09943__A2 (.I(_01526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09945__A1 (.I(_04045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09946__A2 (.I(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09948__A1 (.I(_01536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09948__A2 (.I(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09950__I (.I(_01088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09952__A1 (.I(_04045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09952__B (.I(_04063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09954__B1 (.I(_04065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09954__B2 (.I(_00766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09954__C (.I(_00764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09956__A1 (.I(_04015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09956__A2 (.I(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09958__I (.I(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09960__A1 (.I(_03681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09961__A1 (.I(_01903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09962__A1 (.I(_04037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09964__I (.I(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09966__I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09967__A1 (.I(_04037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09968__A1 (.I(_04077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09970__A1 (.I(_02853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09970__A2 (.I(_00721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09970__B1 (.I(_00889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09970__B2 (.I(_04077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09970__C (.I(_00733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09971__I (.I(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09972__A1 (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09974__A1 (.I(_01912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09976__I (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09977__A1 (.I(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09977__A2 (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09977__B1 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09977__B2 (.I(_01901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09978__A1 (.I(_04087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09978__A2 (.I(_01535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09981__A2 (.I(_04091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09982__A1 (.I(_04077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09982__A2 (.I(_02942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09982__B (.I(_03814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09983__A2 (.I(_04081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09984__A1 (.I(_01913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09984__A2 (.I(_03895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09984__C (.I(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09986__A1 (.I(_04096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09986__A2 (.I(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09987__A1 (.I(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09987__A2 (.I(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09988__A1 (.I(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09988__A2 (.I(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09993__A1 (.I(_02853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09993__C (.I(_04103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09994__A1 (.I(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09994__A2 (.I(_01613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09995__A2 (.I(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__09996__A2 (.I(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10002__A1 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10002__B (.I(_04111_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10002__C (.I(_04112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10003__B (.I(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10004__B (.I(_00598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10008__A1 (.I(_04114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10008__B1 (.I(_04118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10008__B2 (.I(_00866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10009__B (.I(_03865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10010__A1 (.I(_01913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10010__A2 (.I(_03751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10011__I (.I(_00845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10012__A1 (.I(_04077_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10013__A2 (.I(_04121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10014__I (.I(_00826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10015__I (.I(_00718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10016__I (.I(_03766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10017__I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10018__A1 (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10018__A2 (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10019__A1 (.I(_04127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10020__A1 (.I(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10020__B2 (.I(_04127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10020__C (.I(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10021__A1 (.I(_00724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10022__A1 (.I(_01922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10022__A2 (.I(_04126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10023__I (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10024__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10029__A1 (.I(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10029__A2 (.I(_03814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10030__A1 (.I(_04127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10030__A2 (.I(_04038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10031__A1 (.I(_04125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10032__I (.I(_00876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10033__A1 (.I(_01922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10033__A2 (.I(_04017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10036__I (.I(_04096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10037__A1 (.I(_04146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10037__A2 (.I(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10039__A2 (.I(_01713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10040__A1 (.I(_00603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10042__A1 (.I(_04146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10042__A2 (.I(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10044__A2 (.I(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10045__A1 (.I(_00603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10046__C (.I(_03972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10048__I (.I(_00596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10049__B1 (.I(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10051__I (.I(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10052__B2 (.I(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10053__A1 (.I(_01922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10054__A1 (.I(_04127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10056__I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10057__A1 (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10057__A2 (.I(_04096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10061__A1 (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10064__A1 (.I(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10064__A2 (.I(_04172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10065__A1 (.I(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10065__A2 (.I(_02942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10066__I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10068__A1 (.I(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10069__I (.I(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10071__A2 (.I(_04048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10072__A2 (.I(_00631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10073__A1 (.I(_00743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10073__A2 (.I(_04177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10073__C (.I(_00734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10075__A1 (.I(_02185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10075__A2 (.I(_03895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10075__B1 (.I(_04017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10078__A2 (.I(_01701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10079__A2 (.I(_01701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10079__B (.I(_01103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10080__A1 (.I(_04187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10080__A2 (.I(_04188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10081__A1 (.I(_04186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10082__A2 (.I(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10083__A2 (.I(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10084__A1 (.I(_04191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10084__A2 (.I(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10085__A1 (.I(_04186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10087__A1 (.I(_03972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10087__B2 (.I(_04195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10088__A2 (.I(_04177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10088__B2 (.I(_00766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10088__C (.I(_00764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10093__A1 (.I(_00764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10096__A1 (.I(_02185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10098__A1 (.I(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10101__A1 (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10103__A2 (.I(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10108__A1 (.I(_04186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10108__A2 (.I(_04191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10108__A3 (.I(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10109__A1 (.I(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10110__A2 (.I(_04187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10110__A3 (.I(_04188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10112__A1 (.I(_04103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10112__B2 (.I(_04112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10113__I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10114__A1 (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10115__A1 (.I(_04221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10116__A1 (.I(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10116__A2 (.I(_04220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10118__I (.I(_04126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10119__I (.I(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10120__I (.I(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10121__A1 (.I(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10121__B2 (.I(_04221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10121__C (.I(_01231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10123__A1 (.I(_02196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10127__A1 (.I(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10127__A2 (.I(_04234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10128__A1 (.I(_04221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10128__A2 (.I(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10129__A1 (.I(_00719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10130__A1 (.I(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10132__I (.I(_03981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10133__A1 (.I(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10133__B2 (.I(_04240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10134__A1 (.I(_04221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10136__I (.I(_00541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10139__A1 (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10139__A2 (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10140__A1 (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10141__A2 (.I(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10143__I (.I(_04249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10144__I (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10145__I (.I(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10146__B2 (.I(_04251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10147__A1 (.I(_02203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10147__A2 (.I(_04245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10148__A1 (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10150__A1 (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10150__B (.I(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10154__A1 (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10154__B (.I(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10155__A1 (.I(_04244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10156__A1 (.I(_02204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10156__A2 (.I(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10156__B2 (.I(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10156__C (.I(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10157__A2 (.I(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10163__A1 (.I(_04191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10163__A2 (.I(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10166__B (.I(_04272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10167__B (.I(_00636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10168__A1 (.I(_04187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10168__A2 (.I(_04188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10169__B (.I(_04272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10170__B (.I(_03972_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10172__A2 (.I(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10172__B1 (.I(_04278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10172__B2 (.I(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10173__A1 (.I(_00866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10173__A2 (.I(_04268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10174__B (.I(_03865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10175__A1 (.I(_02204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10175__A2 (.I(_03751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10176__I (.I(_00845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10177__A1 (.I(net96));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10177__B (.I(_04283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10178__A2 (.I(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10179__A1 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10179__A2 (.I(_04096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10180__A2 (.I(_04146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10184__A1 (.I(_04289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10187__A1 (.I(_04063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10187__B2 (.I(_04112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10188__A1 (.I(_04251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10189__A1 (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10191__A2 (.I(_04293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10192__A1 (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10192__A2 (.I(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10193__I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10194__A1 (.I(_04289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10194__B2 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10194__C (.I(_01231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10196__A1 (.I(_02209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10200__A1 (.I(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10201__A1 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10201__A2 (.I(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10202__A1 (.I(_00719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10203__A1 (.I(_02210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10205__A1 (.I(_02210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10205__B2 (.I(_04240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10206__A1 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10206__B (.I(_04283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10209__A1 (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10209__A2 (.I(_04146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10212__A1 (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10212__A2 (.I(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10213__A2 (.I(_04317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10214__I (.I(\as2650.addr_buff[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10216__A1 (.I(_04319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10218__A1 (.I(\as2650.addr_buff[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10219__A1 (.I(_04112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10219__B2 (.I(_04063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10220__A1 (.I(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10221__A1 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10223__A1 (.I(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10224__A1 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10224__A2 (.I(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10225__A1 (.I(_04319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10225__A2 (.I(_04020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10226__I (.I(_02515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10228__A1 (.I(_02216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10231__A1 (.I(_04317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10233__A1 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10233__A2 (.I(_04038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10234__A1 (.I(_04125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10235__A1 (.I(_02217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10236__B2 (.I(_00827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10237__A1 (.I(_02217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10237__B2 (.I(_04240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10238__A1 (.I(net95));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10238__B (.I(_04283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10241__A1 (.I(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10244__A1 (.I(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10244__A2 (.I(_00609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10249__A1 (.I(_00638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10249__A2 (.I(_00651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10249__A3 (.I(_00916_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10250__A1 (.I(_00770_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10251__A1 (.I(_00473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10251__A2 (.I(_00544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10253__A1 (.I(_00626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10254__A1 (.I(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10254__A2 (.I(_00885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10255__A1 (.I(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10256__A1 (.I(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10256__A2 (.I(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10256__A3 (.I(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10257__A1 (.I(_03613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10259__A1 (.I(_04346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10260__A2 (.I(_04345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10262__I (.I(_00791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10264__I (.I(_04367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10265__A1 (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10265__A2 (.I(_04368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10266__A1 (.I(_03927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10266__A2 (.I(_00503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10267__A1 (.I(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10269__A1 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10269__A2 (.I(_04372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10269__A3 (.I(_04017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10270__A1 (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10270__A2 (.I(_00592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10270__B (.I(_00654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10270__C (.I(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10271__A1 (.I(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10272__A1 (.I(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10273__A1 (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10273__C (.I(_03689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10274__A1 (.I(_00782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10274__A2 (.I(_00893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10274__A3 (.I(_00726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10276__A1 (.I(_04378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10277__A2 (.I(_00738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10277__A3 (.I(_00491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10277__A4 (.I(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10278__A1 (.I(_00738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10278__A2 (.I(_00708_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10281__A1 (.I(_00679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10281__A3 (.I(_00732_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10281__A4 (.I(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10282__A1 (.I(_00738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10283__A2 (.I(_00695_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10285__A1 (.I(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10285__A2 (.I(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10289__A1 (.I(_02739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10289__A2 (.I(_02932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10290__A1 (.I(_00838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10290__A2 (.I(_00829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10290__A3 (.I(_02506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10291__A3 (.I(_03766_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10292__A1 (.I(_00782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10292__A2 (.I(_00466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10293__B (.I(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10295__A2 (.I(_03719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10295__A4 (.I(_04397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10296__A2 (.I(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10297__I (.I(_00710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10298__A2 (.I(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10299__A2 (.I(_00647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10299__A3 (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10299__B1 (.I(_00721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10301__A1 (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10301__B (.I(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10302__A1 (.I(_00861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10302__A2 (.I(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10303__I (.I(_00805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10304__A1 (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10304__A2 (.I(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10305__A1 (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10305__A4 (.I(_03810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10306__A1 (.I(_03729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10306__A3 (.I(_04407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10307__B (.I(_02548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10308__A1 (.I(net94));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10308__B (.I(_04283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10309__A2 (.I(_04410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10310__I (.I(_03109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10311__A1 (.I(_00829_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10311__A2 (.I(_00709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10312__A1 (.I(_00724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10312__A2 (.I(_00701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10312__B1 (.I(_04413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10312__B2 (.I(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10313__A1 (.I(_00609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10313__A2 (.I(_03723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10314__A1 (.I(_00917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10317__A1 (.I(_00541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10317__A2 (.I(_00800_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10317__A3 (.I(_04418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10318__I (.I(_01033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10319__A1 (.I(_00844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10319__A2 (.I(_00654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10319__C (.I(_04420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10320__A1 (.I(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10322__B2 (.I(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10325__A1 (.I(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10326__A1 (.I(_00627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10326__A2 (.I(_00733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10326__A3 (.I(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10327__A1 (.I(_00536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10327__B (.I(_04424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10328__I (.I(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10329__I (.I(_04430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10330__I (.I(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10332__A1 (.I(_04412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10333__I (.I(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10335__A1 (.I(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10336__A1 (.I(_04272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10337__A1 (.I(_03884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10338__A1 (.I(_04289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10339__A1 (.I(_03951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10340__I (.I(_04319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10341__A1 (.I(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10342__A1 (.I(_04003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10343__I (.I(_01036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10344__A1 (.I(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10344__A2 (.I(_04430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10345__A1 (.I(_03203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10346__I (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10347__I (.I(_01035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10348__I0 (.I(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10348__I1 (.I(_04443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10348__S (.I(_04430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10349__I (.I(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10350__A2 (.I(_04430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10351__A1 (.I(_04038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10352__A2 (.I(_04033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10353__A2 (.I(_02548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10353__C (.I(_03689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10354__I (.I(_00914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10355__A1 (.I(_04447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10355__B (.I(_02537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10355__C (.I(_03689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10357__A1 (.I(_00596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10358__A1 (.I(_00624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10358__A2 (.I(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10358__B1 (.I(_02536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10358__B2 (.I(_02490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10359__A1 (.I(_04378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10362__A1 (.I(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10362__A2 (.I(_00638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10363__A2 (.I(_00756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10363__A3 (.I(_00917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10363__A4 (.I(_03729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10365__A1 (.I(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10365__A2 (.I(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10365__B (.I(_04456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10366__I (.I(_03688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10367__A2 (.I(_04456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10367__B (.I(_04457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10367__C (.I(_04458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10368__A1 (.I(_04443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10368__A2 (.I(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10368__B (.I(_04456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10369__A2 (.I(_04456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10369__B (.I(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10369__C (.I(_04458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10370__A1 (.I(_00792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10370__A2 (.I(_02856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10371__A2 (.I(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10371__B (.I(_04460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10372__A1 (.I(_00902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10372__A2 (.I(_00961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10372__C (.I(_01117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10373__B (.I(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10374__A1 (.I(_00894_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10374__A2 (.I(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10375__I (.I(_04464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10376__I0 (.I(_04461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10376__S (.I(_04465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10378__A1 (.I(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10378__A2 (.I(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10380__A1 (.I(_01850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10380__A2 (.I(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10381__A1 (.I(_04467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10382__I0 (.I(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10382__S (.I(_04465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10384__I (.I(_04464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10385__I (.I(_00792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10386__I (.I(_04473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10387__A1 (.I(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10387__A2 (.I(_03884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10388__A1 (.I(_02067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10388__A2 (.I(_00796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10388__B (.I(_04475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10389__I (.I(_04464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10391__A2 (.I(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10392__A1 (.I(_00794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10392__A2 (.I(_03951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10393__A1 (.I(_02098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10393__A2 (.I(_00796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10395__A2 (.I(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10396__A1 (.I(_00537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10396__A2 (.I(_04003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10397__A1 (.I(_03622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10397__A2 (.I(_00796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10399__A2 (.I(_04483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10401__A1 (.I(_01899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10401__A2 (.I(_00583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10402__A1 (.I(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10402__A2 (.I(_04045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10403__A2 (.I(_04465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10404__A2 (.I(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10405__I (.I(_03927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10406__A1 (.I(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10406__A2 (.I(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10407__A1 (.I(_03625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10407__A2 (.I(_04489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10408__I1 (.I(\as2650.holding_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10408__S (.I(_04464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10411__A1 (.I(_04489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10411__A2 (.I(_00852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10411__B (.I(_04465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10412__B2 (.I(_02345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10413__I (.I(_00838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10414__A1 (.I(_04495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10414__A2 (.I(_00853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10415__B (.I(_00668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10418__A2 (.I(_02857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10418__B (.I(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10419__A2 (.I(_04498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10419__B (.I(_04500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10420__I (.I(_02858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10421__A2 (.I(_04501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10421__B (.I(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10422__A1 (.I(_05725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10422__A2 (.I(_04498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10422__B (.I(_04502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10423__I (.I(_02860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10424__A1 (.I(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10424__B1 (.I(_04498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10426__A1 (.I(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10426__A2 (.I(_00854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10426__B (.I(_00668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10427__A2 (.I(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10427__B (.I(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10428__A1 (.I(_01108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10430__A1 (.I(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10430__B1 (.I(_04498_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10430__B2 (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10432__A1 (.I(_00852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10432__B2 (.I(_01180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10434__A2 (.I(_03736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10435__A1 (.I(_00624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10435__A2 (.I(_00823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10435__A3 (.I(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10436__A1 (.I(_04510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10436__B (.I(_00773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10438__A1 (.I(_02520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10439__A1 (.I(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10440__A1 (.I(_02538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10441__A1 (.I(_04346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10443__A1 (.I(_03613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10444__A2 (.I(_00721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10444__A3 (.I(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10444__A4 (.I(_04418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10445__A1 (.I(_02523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10445__A2 (.I(_04510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10448__A1 (.I(_02504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10448__A2 (.I(_04345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10449__I (.I(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10452__A1 (.I(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10454__I (.I(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10455__I (.I(_00583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10456__A1 (.I(_01836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10456__A2 (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10457__A1 (.I(_00626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10457__A2 (.I(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10458__A2 (.I(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10460__A2 (.I(_04534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10461__A1 (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10462__A1 (.I(_04532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10463__A1 (.I(_00458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10464__A2 (.I(_00458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10465__B2 (.I(_04532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10466__I (.I(_04413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10467__A2 (.I(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10468__A1 (.I(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10468__A2 (.I(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10469__A1 (.I(_04541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10470__A1 (.I(_04412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10470__A2 (.I(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10471__A1 (.I(_04186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10472__B (.I(_00793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10473__A1 (.I(_04530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10473__C (.I(_00740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10474__I (.I(_01231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10475__A1 (.I(_05832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10475__A2 (.I(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10476__A1 (.I(_02856_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10476__B (.I(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10477__A1 (.I(_03768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10478__I (.I(_00512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10479__A1 (.I(_01836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10479__A2 (.I(_04549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10479__B (.I(_04552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10479__C (.I(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10480__A1 (.I(_04244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10482__A1 (.I(_03927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10484__I (.I(_04558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10486__I (.I(_01809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10488__I (.I(_01952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10490__A1 (.I(\as2650.stack[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10490__B1 (.I(_04564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10494__A1 (.I(\as2650.stack[11][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10494__A2 (.I(_04566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10494__B1 (.I(_04568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10494__B2 (.I(\as2650.stack[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10495__A1 (.I(_04560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10497__A1 (.I(\as2650.stack[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10497__A2 (.I(_04566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10497__B1 (.I(_04568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10497__B2 (.I(\as2650.stack[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10500__A2 (.I(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10500__B1 (.I(_04574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10500__B2 (.I(\as2650.stack[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10501__A1 (.I(_04571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10503__A1 (.I(\as2650.stack[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10503__B2 (.I(\as2650.stack[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10504__A1 (.I(\as2650.stack[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10506__A2 (.I(_02837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10507__A2 (.I(_02835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10507__B1 (.I(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10507__B2 (.I(\as2650.stack[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10508__A1 (.I(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10509__B (.I(_01943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10511__A1 (.I(_04559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10511__A2 (.I(_04585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10513__I (.I(_04587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10514__B (.I(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10515__A1 (.I(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10516__A1 (.I(_01791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10518__B1 (.I(_04591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10518__C (.I(_04592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10519__A2 (.I(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10519__C (.I(_04458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10521__I (.I(_04587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10522__I (.I(_01809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10523__I (.I(_01952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10524__A1 (.I(\as2650.stack[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10524__B2 (.I(\as2650.stack[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10525__A1 (.I(\as2650.stack[11][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10525__B2 (.I(\as2650.stack[10][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10527__A1 (.I(\as2650.stack[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10527__B2 (.I(\as2650.stack[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10528__A1 (.I(\as2650.stack[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10528__B2 (.I(\as2650.stack[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10532__A1 (.I(\as2650.stack[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10532__B2 (.I(\as2650.stack[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10534__A1 (.I(\as2650.stack[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10534__B2 (.I(\as2650.stack[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10535__B2 (.I(\as2650.stack[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10537__B (.I(_01942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10538__A1 (.I(_02817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10539__A2 (.I(_04612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10540__I (.I(_04558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10541__A2 (.I(_04594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10541__B (.I(_03754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10542__I (.I(_00473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10543__A2 (.I(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10544__A1 (.I(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10544__A2 (.I(_03821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10545__A1 (.I(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10545__A2 (.I(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10545__B (.I(_00895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10546__A1 (.I(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10547__A1 (.I(_04413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10547__B1 (.I(_04594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10550__A1 (.I(_03809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10551__A1 (.I(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10551__A2 (.I(_04534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10553__A1 (.I(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10553__A2 (.I(_04534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10554__A2 (.I(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10555__A1 (.I(_02549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10556__A1 (.I(_00584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10557__I (.I(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10558__I (.I(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10559__A1 (.I(_01079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10559__A2 (.I(_05832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10560__A2 (.I(_05826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10561__A2 (.I(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10561__B (.I(_04020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10562__A2 (.I(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10563__A1 (.I(_02858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10563__B (.I(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10564__A2 (.I(_04594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10565__A1 (.I(_04632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10567__A1 (.I(_04640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10567__A2 (.I(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10568__A1 (.I(_04367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10570__A1 (.I(_04616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10570__B2 (.I(_04372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10572__A1 (.I(_04591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10572__A2 (.I(_04594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10572__C (.I(_04592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10573__A1 (.I(_03809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10573__A2 (.I(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10573__C (.I(_04458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10574__I (.I(_04591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10576__A2 (.I(_04648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10577__A1 (.I(\as2650.stack[8][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10577__A2 (.I(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10577__B1 (.I(_02962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10577__B2 (.I(\as2650.stack[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10578__A1 (.I(\as2650.stack[11][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10578__A2 (.I(_02951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10578__B1 (.I(_02957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10578__B2 (.I(\as2650.stack[10][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10579__A1 (.I(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10580__A1 (.I(\as2650.stack[15][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10580__B1 (.I(_02957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10581__A2 (.I(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10581__B1 (.I(_02962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10582__A1 (.I(_02950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10584__A2 (.I(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10584__B1 (.I(_02962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10585__A1 (.I(\as2650.stack[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10587__A1 (.I(\as2650.stack[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10587__B2 (.I(\as2650.stack[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10588__A1 (.I(\as2650.stack[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10588__B2 (.I(\as2650.stack[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10589__A1 (.I(_02950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10590__B (.I(_02817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10591__A1 (.I(_01943_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10592__A1 (.I(_02567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10592__A2 (.I(_04664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10593__I (.I(_04558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10595__A2 (.I(_04649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10595__B (.I(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10596__I (.I(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10597__I (.I(_02932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10601__A1 (.I(_04541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10601__A2 (.I(_04672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10601__B1 (.I(_04649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10601__B2 (.I(_04245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10601__C (.I(_04673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10602__A1 (.I(_01866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10602__A2 (.I(_04648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10603__A1 (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10606__A1 (.I(_04530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10610__A1 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10610__A2 (.I(_05819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10611__A1 (.I(_01214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10611__A2 (.I(_05826_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10612__A2 (.I(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10614__B (.I(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10615__A1 (.I(_02859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10616__A1 (.I(_04686_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10616__A2 (.I(_04687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10617__A1 (.I(_04682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10619__A1 (.I(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10620__A2 (.I(_04672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10621__A1 (.I(_03754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10622__A1 (.I(_04616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10622__B2 (.I(_00741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10627__A2 (.I(_04649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10628__I (.I(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10630__A1 (.I(_01868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10630__B (.I(_04702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10632__I (.I(_04413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10633__A1 (.I(_03921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10633__A2 (.I(_00604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10634__A1 (.I(_02942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10635__A2 (.I(_04706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10636__A1 (.I(_01866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10636__A2 (.I(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10636__A3 (.I(_01834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10637__A1 (.I(_01877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10638__A1 (.I(_03951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10638__A2 (.I(_00743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10640__A1 (.I(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10640__A2 (.I(_00928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10640__B (.I(_00748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10641__A2 (.I(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10641__C (.I(_04368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10642__I (.I(_00715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10643__A1 (.I(_03921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10645__I (.I(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10646__I (.I(_04473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10647__A2 (.I(_04717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10647__B (.I(_04718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10648__A1 (.I(_00462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10650__A2 (.I(_04717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10651__A1 (.I(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10651__A2 (.I(_04706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10651__C (.I(_00543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10652__A2 (.I(_05811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10653__A1 (.I(_01264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10653__A2 (.I(_05819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10656__A1 (.I(_04724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10657__A1 (.I(_04724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10658__A1 (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10658__A2 (.I(_04729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10659__A1 (.I(_02863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10659__A2 (.I(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10660__A1 (.I(_04728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10660__C (.I(_04682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10661__A2 (.I(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10661__C (.I(_04372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10662__A1 (.I(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10665__A1 (.I(\as2650.stack[8][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10665__A2 (.I(_04735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10665__B1 (.I(_04736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10665__B2 (.I(\as2650.stack[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10666__A1 (.I(\as2650.stack[11][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10666__A2 (.I(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10666__B1 (.I(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10666__B2 (.I(\as2650.stack[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10667__A1 (.I(_04560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10669__A1 (.I(\as2650.stack[15][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10669__A2 (.I(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10669__B1 (.I(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10670__A2 (.I(_04735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10670__B1 (.I(_04736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10670__B2 (.I(\as2650.stack[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10671__A1 (.I(_01970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10673__A1 (.I(\as2650.stack[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10673__A2 (.I(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10673__B1 (.I(_04574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10674__A2 (.I(_02824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10674__B1 (.I(_04568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10674__B2 (.I(\as2650.stack[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10676__A2 (.I(_02824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10676__B1 (.I(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10676__B2 (.I(\as2650.stack[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10677__A2 (.I(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10677__B1 (.I(_04574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10677__B2 (.I(\as2650.stack[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10678__A1 (.I(_04571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10679__B (.I(_02946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10681__A2 (.I(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10682__A1 (.I(_02567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10682__A2 (.I(_04717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10682__C (.I(_00877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10684__A2 (.I(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10685__I (.I(_00507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10686__A1 (.I(_01877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10686__A2 (.I(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10686__C (.I(_04757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10688__A1 (.I(_03920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10689__A1 (.I(_04014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10690__A1 (.I(_04015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10691__A1 (.I(_00462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10692__A1 (.I(_01877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10693__A1 (.I(_04014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10694__A1 (.I(_00888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10694__A2 (.I(_04764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10694__B (.I(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10695__A1 (.I(_04015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10696__A1 (.I(_00604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10696__A2 (.I(_04026_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10697__A1 (.I(_04319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10698__A1 (.I(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10698__B (.I(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10699__B (.I(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10700__A2 (.I(_04764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10700__B1 (.I(_04767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10702__I (.I(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10703__A1 (.I(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10703__A2 (.I(_04048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10704__A2 (.I(_05801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10705__A1 (.I(_02862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10705__A2 (.I(_05811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10706__A1 (.I(_04724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10709__A1 (.I(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10710__A2 (.I(_04780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10710__B (.I(_04773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10711__A1 (.I(_04773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10711__A2 (.I(_04764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10712__A1 (.I(_01889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10713__A1 (.I(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10714__A1 (.I(_00537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10714__A2 (.I(_04767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10714__C (.I(_04244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10715__A1 (.I(_00514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10715__C (.I(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10716__A1 (.I(\as2650.stack[8][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10716__B1 (.I(_04564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10716__B2 (.I(\as2650.stack[9][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10717__A1 (.I(\as2650.stack[11][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10717__A2 (.I(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10717__B1 (.I(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10718__A1 (.I(_04560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10719__A1 (.I(\as2650.stack[15][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10719__A2 (.I(_04566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10719__B1 (.I(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10720__A1 (.I(\as2650.stack[12][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10720__B1 (.I(_04564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10720__B2 (.I(\as2650.stack[13][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10721__A1 (.I(_04571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10723__A1 (.I(\as2650.stack[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10724__A1 (.I(\as2650.stack[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10724__B1 (.I(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10727__A2 (.I(_02835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10727__B1 (.I(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10727__B2 (.I(\as2650.stack[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10728__A1 (.I(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10729__B (.I(_02946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10731__A2 (.I(_04801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10732__A1 (.I(_02567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10732__C (.I(_00877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10734__A2 (.I(_04764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10735__I (.I(_03688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10736__A1 (.I(_01889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10739__I (.I(_04808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10740__A1 (.I(\as2650.stack[8][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10740__A2 (.I(_04735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10740__B1 (.I(_04736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10740__B2 (.I(\as2650.stack[9][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10741__A1 (.I(\as2650.stack[11][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10741__A2 (.I(_01980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10741__B1 (.I(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10742__A1 (.I(_01949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10743__A1 (.I(\as2650.stack[15][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10743__A2 (.I(_01980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10743__B1 (.I(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10744__A2 (.I(_04735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10744__B1 (.I(_04736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10745__A1 (.I(_01970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10747__A1 (.I(\as2650.stack[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10747__B1 (.I(_04564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10748__A1 (.I(\as2650.stack[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10748__A2 (.I(_04566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10748__B1 (.I(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10749__A1 (.I(_04560_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10750__A1 (.I(\as2650.stack[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10750__A2 (.I(_02824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10750__B1 (.I(_04568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10751__A2 (.I(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10751__B1 (.I(_04574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10751__B2 (.I(\as2650.stack[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10752__A1 (.I(_04571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10753__B (.I(_02946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10754__A1 (.I(_01944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10755__A2 (.I(_04824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10756__I (.I(_00876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10759__A1 (.I(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10759__A2 (.I(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10760__A1 (.I(_01535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10760__A2 (.I(_05789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10761__A2 (.I(_05801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10764__B (.I(_00787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10766__B (.I(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10767__A1 (.I(_04549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10767__A2 (.I(_04808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10767__B (.I(_04836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10769__A2 (.I(_04808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10771__A1 (.I(_00602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10771__A2 (.I(_04042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10772__A1 (.I(_01903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10772__A2 (.I(_00849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10772__B (.I(_04841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10773__A1 (.I(_01036_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10774__A1 (.I(_03203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10775__A2 (.I(_04808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10775__B1 (.I(_04844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10775__B2 (.I(_00895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10775__C (.I(_00792_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10776__A1 (.I(_00859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10777__A1 (.I(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10777__A2 (.I(_04840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10778__C (.I(_00853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10779__A1 (.I(_00536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10780__A1 (.I(_04718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10781__A1 (.I(_03754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10782__B (.I(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10783__A1 (.I(_03680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10783__C (.I(_00777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10784__I (.I(_01791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10786__I (.I(_02521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10789__A1 (.I(_04087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10790__I (.I(_01912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10794__I (.I(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10795__A1 (.I(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10795__A2 (.I(_05857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10796__A2 (.I(_05789_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10799__B (.I(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10800__A1 (.I(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10800__A2 (.I(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10802__A1 (.I(_01912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10802__A2 (.I(_01901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10803__A1 (.I(_04860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10805__A2 (.I(_04873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10806__A1 (.I(_04863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10806__A2 (.I(_04870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10807__A1 (.I(_01901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10807__A2 (.I(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10808__A1 (.I(_04860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10810__A2 (.I(_04873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10810__C (.I(_04473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10811__A1 (.I(_00849_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10811__A2 (.I(_04091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10812__A1 (.I(_01913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10813__A1 (.I(_04443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10814__A1 (.I(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10814__A2 (.I(_00699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10815__A1 (.I(_04882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10816__I (.I(_00791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10817__A2 (.I(_04862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10817__B2 (.I(_00710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10817__C (.I(_04885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10818__A1 (.I(_00860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10818__B (.I(_04886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10819__A1 (.I(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10820__C (.I(_00853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10821__I (.I(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10822__A2 (.I(_04862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10823__C (.I(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10824__A1 (.I(_00834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10825__A2 (.I(_04873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10826__A2 (.I(_02846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10827__A1 (.I(_00827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10828__A1 (.I(_03680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10828__A2 (.I(_04862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10828__C (.I(_00777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10829__A1 (.I(\as2650.ivec[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10829__B2 (.I(_04862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10830__A1 (.I(_04860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10832__A1 (.I(_04899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10833__I (.I(_04900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10834__A1 (.I(_04899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10834__A2 (.I(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10835__A1 (.I(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10836__A1 (.I(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10836__A2 (.I(_04020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10837__A1 (.I(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10838__A2 (.I(_04900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10838__B2 (.I(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10838__C (.I(_00793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10839__A1 (.I(_00860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10841__A1 (.I(_04860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10842__A1 (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10843__A1 (.I(_00888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10843__A2 (.I(_04900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10845__B (.I(_00715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10846__A1 (.I(_04530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10847__A1 (.I(_04368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10847__A2 (.I(_04900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10847__C (.I(_04125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10848__A1 (.I(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10849__A1 (.I(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10849__A2 (.I(_05857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10850__A1 (.I(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10850__A2 (.I(_05778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10851__A2 (.I(_04918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10852__B (.I(_04549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10853__A1 (.I(_04773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10853__A2 (.I(_04901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10853__B (.I(_04920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10854__A1 (.I(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10855__A2 (.I(_04901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10856__A2 (.I(_02966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10857__B (.I(_00827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10858__A1 (.I(_03680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10858__A2 (.I(_04901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10858__C (.I(_03865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10859__A1 (.I(\as2650.ivec[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10859__B2 (.I(_04901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10859__C (.I(_04592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10860__A1 (.I(_04899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10861__I (.I(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10862__I (.I(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10863__A1 (.I(_04899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10865__I (.I(_04931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10868__A2 (.I(_04932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10869__A2 (.I(_04172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10872__A1 (.I(_04412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10873__A1 (.I(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10873__A2 (.I(_04939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10874__A2 (.I(_04931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10874__B2 (.I(_00860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10875__A1 (.I(_04616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10876__A1 (.I(_02910_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10876__A2 (.I(_05778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10877__A2 (.I(_05778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10879__A1 (.I(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10879__A2 (.I(_04945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10881__A1 (.I(_04632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10881__A2 (.I(_04932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10882__A1 (.I(_04773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10882__A2 (.I(_04947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10882__C (.I(_04372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10883__A2 (.I(_04931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10883__B (.I(_00718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10884__A1 (.I(_00794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10885__A1 (.I(_04929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10885__A2 (.I(_04942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10885__A4 (.I(_04951_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10886__A2 (.I(_04931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10887__A2 (.I(_01990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10888__A1 (.I(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10888__A2 (.I(_04932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10888__B2 (.I(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10888__C (.I(_02547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10890__A1 (.I(_03736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10890__A2 (.I(_04932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10891__A2 (.I(_03736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10891__C (.I(_03981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10893__A1 (.I(_02185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10894__A1 (.I(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10898__A3 (.I(_00699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10898__A4 (.I(_04945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10899__A1 (.I(_04682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10899__A2 (.I(_04964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10900__A2 (.I(_04962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10900__B1 (.I(_04963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10902__B (.I(_02196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10903__I (.I(_04962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10904__A2 (.I(_04969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10905__A1 (.I(_00888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10906__A1 (.I(_02196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10906__A2 (.I(_00603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10907__A1 (.I(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10907__A2 (.I(_04234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10907__C (.I(_04541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10908__A1 (.I(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10909__A1 (.I(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10910__A2 (.I(_04962_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10910__C (.I(_04367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10911__A1 (.I(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10912__I (.I(_02559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10913__A2 (.I(_04234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10913__C (.I(_03858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10914__A1 (.I(_04978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10914__A2 (.I(_04969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10915__B2 (.I(_00719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10915__C (.I(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10916__A1 (.I(_00741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10917__A1 (.I(_00861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10917__A2 (.I(_04559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10919__A1 (.I(_02042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10919__A2 (.I(_03657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10919__B1 (.I(_04969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10919__C (.I(_04984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10920__B2 (.I(_04969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10921__A1 (.I(_04982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10922__A1 (.I(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10923__A1 (.I(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10925__A1 (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10927__A1 (.I(_02203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10929__A1 (.I(_04272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10931__A2 (.I(_04991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10931__B1 (.I(_04993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10932__I (.I(_04991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10935__A1 (.I(_00462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10935__A2 (.I(_04997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10935__C (.I(_04718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10936__A1 (.I(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10937__A2 (.I(_04964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10938__A2 (.I(_04964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10939__A1 (.I(_04549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10940__A1 (.I(_04632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10940__A2 (.I(_04991_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10941__A1 (.I(_00584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10941__A2 (.I(_04993_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10942__A1 (.I(_04978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10942__A2 (.I(_04997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10943__A1 (.I(_00514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10943__C (.I(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10944__A1 (.I(_04616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10945__A1 (.I(_02065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10945__A2 (.I(_03657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10945__B2 (.I(_04997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10945__C (.I(_04984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10946__B2 (.I(_04997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10947__A1 (.I(_05009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10948__A1 (.I(_02204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10949__A1 (.I(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10952__I (.I(_05015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10953__A1 (.I(_02209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10953__A2 (.I(_00850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10955__A1 (.I(_04978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10956__A1 (.I(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10956__A2 (.I(_05016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10956__C (.I(_04244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10957__A1 (.I(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10958__A1 (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10959__A1 (.I(_02203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10959__B (.I(_02209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10961__I0 (.I(_05016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10963__A1 (.I(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10964__A1 (.I(_04245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10964__A2 (.I(_05015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10964__B2 (.I(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10965__A1 (.I(_04368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10966__A1 (.I(_04249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10966__A2 (.I(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10966__A3 (.I(_04964_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10967__A1 (.I(_04289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10967__B (.I(_04863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10968__A2 (.I(_05016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10968__C (.I(_00830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10969__A1 (.I(_00514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10970__A2 (.I(_05015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10971__A2 (.I(_02095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10971__B (.I(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10972__C (.I(_03681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10973__A1 (.I(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10973__A2 (.I(_05016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10973__B (.I(_04033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10974__B2 (.I(_05015_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10975__A1 (.I(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10977__A1 (.I(_02210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10977__B (.I(_04702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10979__I (.I(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10983__I0 (.I(_02216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10984__I0 (.I(_05045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10984__I1 (.I(_05046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10984__S (.I(_04978_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10985__A1 (.I(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10986__A1 (.I(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10987__A1 (.I(_04632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10987__A2 (.I(_05045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10987__B (.I(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10988__A1 (.I(_02216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10991__C (.I(_04640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10992__A1 (.I(\as2650.addr_buff[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10992__A2 (.I(_00723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10993__B (.I(_04885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10994__A1 (.I(_04126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10994__B1 (.I(_05046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10994__B2 (.I(_00859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10994__C (.I(_05056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10996__C (.I(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10997__A1 (.I(_00543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10997__C (.I(_00861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10998__A1 (.I(_02118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10998__A2 (.I(_03657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10998__B2 (.I(_05045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10999__A1 (.I(\as2650.ivec[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__10999__B2 (.I(_05045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11001__A1 (.I(_02217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11002__A1 (.I(_05042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11003__I (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11006__A1 (.I(_02224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11007__A1 (.I(_04559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11007__A2 (.I(_05068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11008__A2 (.I(_02144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11009__A1 (.I(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11009__B2 (.I(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11010__A1 (.I(_04863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11010__B (.I(_00740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11011__A1 (.I(_02224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11012__A1 (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11014__A2 (.I(_05068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11014__C (.I(_04640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11015__A1 (.I(_02224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11015__A2 (.I(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11016__A2 (.I(_00787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11017__A1 (.I(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11017__B (.I(_00535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11018__A1 (.I(_04126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11018__A2 (.I(_05068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11018__B2 (.I(_00859_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11019__A1 (.I(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11020__A1 (.I(_05071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11020__C (.I(_04125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11021__A1 (.I(_04530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11022__C (.I(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11023__A1 (.I(_00834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11025__A1 (.I(_04591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11025__C (.I(_04592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11026__I (.I(_03688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11027__A2 (.I(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11027__C (.I(_05088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11029__A1 (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11032__A2 (.I(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11032__B (.I(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11034__A1 (.I(_02231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11035__A1 (.I(_04245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11036__A1 (.I(_02231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11036__A2 (.I(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11037__A1 (.I(_04443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11037__B2 (.I(_04541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11037__C (.I(_04367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11038__A1 (.I(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11038__C (.I(_00740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11039__A1 (.I(_04863_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11040__A1 (.I(_04682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11040__A2 (.I(_04882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11041__A1 (.I(_00543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11042__S (.I(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11043__A1 (.I(_00854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11043__B (.I(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11046__A1 (.I(_02231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11046__B (.I(_04702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11048__A1 (.I(_00475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11048__A2 (.I(_00895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11048__B (.I(_00630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11049__A1 (.I(_00769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11049__C (.I(_00615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11050__A1 (.I(_00638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11050__A2 (.I(_00917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11052__A1 (.I(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11053__A1 (.I(_01118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11053__A2 (.I(_02559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11053__B (.I(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11054__A1 (.I(_00995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11054__B1 (.I(_02761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11055__A1 (.I(_00902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11056__A1 (.I(_00884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11057__B (.I(_04495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11059__A1 (.I(_00675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11059__A2 (.I(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11059__A3 (.I(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11061__A1 (.I(_02739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11061__A2 (.I(_00503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11061__A3 (.I(_00893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11063__A2 (.I(_00893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11063__A3 (.I(_00982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11064__A1 (.I(_00523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11064__B3 (.I(_00680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11066__A2 (.I(_00902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11067__A1 (.I(_00837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11067__A2 (.I(_03723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11069__A1 (.I(_02536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11069__A3 (.I(_05128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11071__A1 (.I(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11074__A1 (.I(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11074__A2 (.I(_01094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11075__I (.I(_00636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11076__I (.I(_00805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11077__A1 (.I(_05135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11077__A2 (.I(_01051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11078__A1 (.I(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11078__A2 (.I(net82));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11078__C (.I(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11079__I (.I(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11080__I (.I(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11081__I (.I(_00982_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11083__A2 (.I(_04585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11084__I (.I(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11085__I (.I(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11086__A1 (.I(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11087__A1 (.I(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11087__B (.I(_01928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11089__I (.I(_00685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11090__A1 (.I(_01146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11091__I (.I(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11094__A1 (.I(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11094__B1 (.I(_05150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11094__C (.I(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11095__A1 (.I(_02857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11095__B (.I(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11097__A1 (.I(_01225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11098__A1 (.I(_00914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11099__A1 (.I(_00455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11099__A2 (.I(_04929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11102__A1 (.I(_01822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11104__A1 (.I(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11106__I (.I(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11107__A1 (.I(\as2650.stack[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11107__A2 (.I(_05166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11108__I (.I(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11109__I (.I(_02131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11110__I (.I(_02132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11111__A1 (.I(\as2650.stack[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11111__B1 (.I(_05169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11111__B2 (.I(\as2650.stack[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11111__C2 (.I(_05170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11112__A1 (.I(_05165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11116__A1 (.I(\as2650.stack[11][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11116__A2 (.I(_05175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11117__I (.I(_02137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11118__A2 (.I(_05177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11118__B1 (.I(_05170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11118__B2 (.I(\as2650.stack[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11118__C1 (.I(\as2650.stack[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11119__A1 (.I(_05174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11121__I (.I(_02083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11122__A1 (.I(\as2650.stack[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11122__A2 (.I(_05181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11123__B1 (.I(_02004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11123__C2 (.I(_02005_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11124__A1 (.I(_05165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11126__I (.I(_02132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11127__A1 (.I(\as2650.stack[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11127__A2 (.I(_05186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11128__B1 (.I(_05169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11128__B2 (.I(\as2650.stack[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11129__A1 (.I(\as2650.stack[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11129__A2 (.I(_05177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11130__A1 (.I(_05185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11132__B (.I(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11133__A1 (.I(_05163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11134__I (.I(_04495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11135__I (.I(_05194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11136__A1 (.I(_05138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11136__A2 (.I(_05159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11136__B1 (.I(_05193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11136__B2 (.I(_05195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11137__A1 (.I(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11137__C (.I(_05088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11138__I (.I(_04420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11139__I (.I(_04063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11140__A1 (.I(_04103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11141__A2 (.I(_01199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11141__C (.I(_04420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11142__A2 (.I(net81));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11142__B (.I(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11143__I0 (.I(_01845_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11143__I1 (.I(_01822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11145__A2 (.I(_04612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11146__C (.I(_02749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11147__A1 (.I(_01237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11147__C (.I(_00685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11148__A1 (.I(_00830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11148__A2 (.I(_05835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11150__A1 (.I(_01212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11150__A2 (.I(_00963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11151__A1 (.I(_04501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11151__B (.I(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11152__A1 (.I(_00454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11152__A2 (.I(_00467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11152__B1 (.I(_03866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11152__B2 (.I(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11153__A1 (.I(_05201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11153__B (.I(_04447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11155__I (.I(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11158__I (.I(_02008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11159__A1 (.I(\as2650.stack[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11159__A2 (.I(_05217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11160__I (.I(_02087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11161__I (.I(_02089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11162__I (.I(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11163__A1 (.I(\as2650.stack[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11163__A2 (.I(_05219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11163__B1 (.I(_05220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11163__B2 (.I(\as2650.stack[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11163__C1 (.I(\as2650.stack[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11163__C2 (.I(_05221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11164__A1 (.I(_05216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11166__I (.I(_02021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11167__A1 (.I(\as2650.stack[11][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11167__A2 (.I(_05225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11168__I (.I(_02126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11169__A1 (.I(\as2650.stack[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11169__A2 (.I(_05227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11169__B1 (.I(_05221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11169__B2 (.I(\as2650.stack[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11169__C1 (.I(\as2650.stack[10][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11169__C2 (.I(_05219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11172__I (.I(_02025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11173__A1 (.I(\as2650.stack[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11173__A2 (.I(_05231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11174__I (.I(_02129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11175__I (.I(_02131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11176__A1 (.I(\as2650.stack[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11176__A2 (.I(_05233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11176__B1 (.I(_05234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11176__B2 (.I(\as2650.stack[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11176__C2 (.I(_05186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11177__A1 (.I(_05216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11178__I (.I(_02061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11179__A2 (.I(_05237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11180__I (.I(_02129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11181__A1 (.I(\as2650.stack[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11181__A2 (.I(_05239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11181__B1 (.I(_05234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11181__B2 (.I(\as2650.stack[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11182__A2 (.I(_05166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11183__A1 (.I(_05185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11185__B (.I(_05243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11186__I (.I(_00914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11187__B (.I(_05244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11187__C (.I(_05245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11188__A2 (.I(_05246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11189__I (.I(_00507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11190__A1 (.I(_01851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11190__B1 (.I(_05212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11191__A1 (.I(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11191__A2 (.I(_01254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11192__A2 (.I(_01260_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11193__A1 (.I(_00806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11193__A2 (.I(net80));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11193__B (.I(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11194__I (.I(_00434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11195__I (.I(_02749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11196__I0 (.I(_01861_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11196__I1 (.I(_01936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11197__A2 (.I(_04664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11199__A1 (.I(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11199__A2 (.I(_05253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11200__A1 (.I(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11201__A1 (.I(_05252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11203__A1 (.I(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11204__I (.I(_00913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11205__A1 (.I(_00441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11205__A2 (.I(_00907_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11205__B (.I(_05262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11206__A1 (.I(_00450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11206__A2 (.I(_03837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11206__B1 (.I(_03810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11209__A2 (.I(_05266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11210__I (.I(_02059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11211__I (.I(_02061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11212__A2 (.I(_05268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11212__B1 (.I(_05175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11212__B2 (.I(\as2650.stack[15][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11212__C2 (.I(_05269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11213__A1 (.I(_05265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11215__I (.I(_02004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11216__A1 (.I(\as2650.stack[11][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11216__A2 (.I(_05273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11217__I (.I(_02080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11218__I (.I(_02059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11219__A1 (.I(\as2650.stack[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11219__A2 (.I(_05181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11219__B1 (.I(_05275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11219__B2 (.I(\as2650.stack[8][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11219__C1 (.I(\as2650.stack[10][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11219__C2 (.I(_05276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11220__A1 (.I(_05272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11223__A1 (.I(\as2650.stack[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11223__A2 (.I(_05266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11224__I (.I(_02082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11225__A1 (.I(\as2650.stack[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11225__A2 (.I(_05282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11225__B1 (.I(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11225__B2 (.I(\as2650.stack[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11225__C1 (.I(\as2650.stack[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11226__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11227__A2 (.I(_05237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11228__I (.I(_02082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11229__I (.I(_01814_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11230__A2 (.I(_05286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11230__B1 (.I(_05287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11230__B2 (.I(\as2650.stack[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11231__A2 (.I(_05231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11232__A1 (.I(_05174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11233__B (.I(_05243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11234__B (.I(_05291_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11235__I (.I(_05194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11236__A1 (.I(_05251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11236__A2 (.I(_05264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11236__B1 (.I(_05292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11237__A1 (.I(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11239__A1 (.I(_02067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11239__B (.I(_05296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11241__A1 (.I(_04195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11241__A2 (.I(_03958_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11242__A1 (.I(_05135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11242__A2 (.I(_01343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11243__A1 (.I(_00806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11243__A2 (.I(_01373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11243__B (.I(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11245__I0 (.I(_01872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11245__I1 (.I(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11245__S (.I(_00939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11246__A2 (.I(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11247__C (.I(_05253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11248__A1 (.I(_01391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11248__B (.I(_05304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11249__A1 (.I(_00441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11250__A1 (.I(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11250__C (.I(_02902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11251__A1 (.I(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11251__A2 (.I(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11251__B (.I(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11252__A1 (.I(_05252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11252__A2 (.I(_03866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11252__B (.I(_05262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11253__A1 (.I(_00452_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11253__A2 (.I(_03837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11254__A1 (.I(\as2650.stack[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11254__A2 (.I(_05266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11255__A2 (.I(_05268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11255__B1 (.I(_05287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11255__B2 (.I(\as2650.stack[15][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11255__C2 (.I(_05269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11256__A1 (.I(_05265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11257__A1 (.I(\as2650.stack[11][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11257__A2 (.I(_05273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11258__A1 (.I(\as2650.stack[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11258__A2 (.I(_05227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11258__B1 (.I(_05275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11258__B2 (.I(\as2650.stack[8][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11258__C1 (.I(\as2650.stack[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11258__C2 (.I(_05268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11259__A1 (.I(_05272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11261__A1 (.I(\as2650.stack[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11261__A2 (.I(_05217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11262__A1 (.I(\as2650.stack[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11262__A2 (.I(_05282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11262__B1 (.I(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11263__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11264__A1 (.I(\as2650.stack[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11264__A2 (.I(_05237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11265__A1 (.I(\as2650.stack[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11265__A2 (.I(_05286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11265__B1 (.I(_05287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11266__A2 (.I(_05166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11267__A1 (.I(_05174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11268__B (.I(_05243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11269__B (.I(_05325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11270__A1 (.I(_05300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11270__A2 (.I(_05310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11270__B1 (.I(_05326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11271__A1 (.I(_02098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11271__B (.I(_05296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11273__A1 (.I(_05135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11273__A2 (.I(_01413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11274__A2 (.I(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11274__B (.I(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11275__A1 (.I(_00806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11275__A2 (.I(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11275__C (.I(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11276__A1 (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11276__A2 (.I(_00939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11277__A1 (.I(_01008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11279__A2 (.I(_04801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11280__A1 (.I(_01724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11280__B (.I(_00685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11281__A1 (.I(_05253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11282__A1 (.I(_05252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11283__A1 (.I(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11283__C (.I(_02902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11284__A1 (.I(_02850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11284__B (.I(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11285__I (.I(_05805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11286__A1 (.I(_05341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11286__A2 (.I(_03866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11286__B (.I(_05262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11287__A1 (.I(_00437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11287__A2 (.I(_03837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11288__A1 (.I(\as2650.stack[13][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11288__A2 (.I(_05266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11289__A2 (.I(_05286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11289__B1 (.I(_05287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11289__B2 (.I(\as2650.stack[15][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11289__C1 (.I(\as2650.stack[12][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11289__C2 (.I(_05275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11290__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11291__A1 (.I(\as2650.stack[11][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11291__A2 (.I(_05273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11292__A1 (.I(\as2650.stack[9][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11292__A2 (.I(_05227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11292__B1 (.I(_05275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11292__B2 (.I(\as2650.stack[8][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11292__C2 (.I(_05268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11295__A1 (.I(\as2650.stack[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11295__A2 (.I(_05217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11296__A2 (.I(_05282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11296__B1 (.I(_05220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11297__A1 (.I(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11298__A1 (.I(\as2650.stack[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11298__A2 (.I(_05237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11299__A2 (.I(_05286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11299__B1 (.I(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11299__B2 (.I(\as2650.stack[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11300__A2 (.I(_05166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11301__A1 (.I(_05174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11302__B (.I(_05243_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11304__A1 (.I(_05331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11304__A2 (.I(_05343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11304__B1 (.I(_05359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11305__A1 (.I(_03622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11305__B (.I(_05296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11307__A1 (.I(_04195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11307__A2 (.I(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11308__A1 (.I(_04103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11308__A2 (.I(_01526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11309__B (.I(_04420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11310__A2 (.I(_01514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11311__A1 (.I(_05341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11313__A1 (.I(_02484_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11314__A2 (.I(_04824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11315__C (.I(_05253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11316__A1 (.I(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11316__A2 (.I(_00984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11316__B (.I(_05370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11318__A1 (.I(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11320__A1 (.I(_02554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11320__C (.I(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11321__A1 (.I(_00428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11321__A2 (.I(_04929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11321__B2 (.I(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11322__A1 (.I(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11323__A1 (.I(_04447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11323__A2 (.I(_05377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11324__A2 (.I(_05217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11325__A2 (.I(_05239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11325__B1 (.I(_05220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11325__B2 (.I(\as2650.stack[15][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11325__C2 (.I(_05221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11326__A1 (.I(_05216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11327__A1 (.I(\as2650.stack[11][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11327__A2 (.I(_05225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11328__A1 (.I(\as2650.stack[9][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11328__A2 (.I(_05177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11328__B1 (.I(_05186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11328__B2 (.I(\as2650.stack[8][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11328__C2 (.I(_05219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11331__A1 (.I(\as2650.stack[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11331__A2 (.I(_05231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11332__A2 (.I(_05233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11332__B1 (.I(_05169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11332__B2 (.I(\as2650.stack[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11332__C2 (.I(_05170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11333__A1 (.I(_05165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11334__A1 (.I(\as2650.stack[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11334__A2 (.I(_05269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11335__A2 (.I(_05239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11335__B1 (.I(_05234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11335__B2 (.I(\as2650.stack[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11336__A2 (.I(_05181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11337__A1 (.I(_05185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11338__B (.I(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11339__A1 (.I(_05163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11339__C (.I(_05245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11341__A1 (.I(_01900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11342__I (.I(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11343__A1 (.I(_05135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11343__A2 (.I(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11344__A2 (.I(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11346__A1 (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11347__A1 (.I(_05735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11347__A2 (.I(_00939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11348__A1 (.I(_01928_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11349__A1 (.I(_01929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11350__A1 (.I(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11351__A1 (.I(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11352__A1 (.I(_02896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11352__C (.I(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11353__A1 (.I(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11353__B (.I(_03653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11354__I (.I(_04495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11355__A1 (.I(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11355__C (.I(_05408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11356__A1 (.I(_00424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11356__A2 (.I(_00467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11356__B1 (.I(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11357__I (.I(_02013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11358__A1 (.I(\as2650.stack[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11358__A2 (.I(_05411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11359__A1 (.I(\as2650.stack[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11359__A2 (.I(_05239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11359__B1 (.I(_05220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11359__B2 (.I(\as2650.stack[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11359__C1 (.I(\as2650.stack[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11359__C2 (.I(_05221_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11360__A1 (.I(_05216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11361__A1 (.I(\as2650.stack[11][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11361__A2 (.I(_05225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11362__A1 (.I(\as2650.stack[9][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11362__A2 (.I(_05177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11362__B1 (.I(_05186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11362__B2 (.I(\as2650.stack[8][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11362__C1 (.I(\as2650.stack[10][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11362__C2 (.I(_05219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11365__A1 (.I(\as2650.stack[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11365__A2 (.I(_05231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11366__A2 (.I(_05233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11366__B1 (.I(_05169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11366__B2 (.I(\as2650.stack[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11366__C2 (.I(_05170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11367__A1 (.I(_05165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11368__A2 (.I(_05269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11369__A2 (.I(_05233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11369__B1 (.I(_05234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11369__B2 (.I(\as2650.stack[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11370__A2 (.I(_05181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11371__A1 (.I(_05185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11372__B (.I(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11373__A1 (.I(_05163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11373__C (.I(_05245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11375__A1 (.I(_03625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11375__B1 (.I(_05410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11376__A1 (.I(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11376__A2 (.I(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11377__A1 (.I(_04195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11377__A2 (.I(_01713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11379__A1 (.I(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11379__A2 (.I(_03228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11379__B (.I(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11380__A1 (.I(_00421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11380__A2 (.I(_04929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11381__A1 (.I(_05727_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11382__A1 (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11383__A2 (.I(_02966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11385__A1 (.I(_03486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11389__A1 (.I(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11389__B1 (.I(_03810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11389__C (.I(_05194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11391__A2 (.I(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11392__A1 (.I(\as2650.stack[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11392__A2 (.I(_05273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11393__I (.I(_02016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11394__A2 (.I(_05411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11394__B1 (.I(_05446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11394__C1 (.I(\as2650.stack[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11394__C2 (.I(_05276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11395__A1 (.I(_05272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11396__A1 (.I(\as2650.stack[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11396__A2 (.I(_05446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11397__A1 (.I(\as2650.stack[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11397__A2 (.I(_05276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11397__B1 (.I(_05175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11397__B2 (.I(\as2650.stack[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11397__C1 (.I(\as2650.stack[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11397__C2 (.I(_05411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11398__A1 (.I(_05265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11400__A2 (.I(_02399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11401__A2 (.I(_05411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11401__B1 (.I(_05446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11401__C1 (.I(\as2650.stack[15][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11401__C2 (.I(_05225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11402__A1 (.I(_05265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11403__A1 (.I(\as2650.stack[9][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11403__A2 (.I(_03027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11404__A2 (.I(_05276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11404__B1 (.I(_05175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11404__B2 (.I(\as2650.stack[11][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11404__C2 (.I(_05446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11405__A1 (.I(_05272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11406__A1 (.I(_05163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11407__A1 (.I(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11408__A1 (.I(_05443_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11409__A1 (.I(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11409__B (.I(_05296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11411__A1 (.I(_04412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11411__A2 (.I(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11412__A1 (.I(_02173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11412__A2 (.I(_02857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11412__B (.I(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11413__A1 (.I(_01054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11413__A2 (.I(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11413__A3 (.I(_00974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11414__A1 (.I(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11414__A2 (.I(_00974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11415__B (.I(_05408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11416__A1 (.I(_00875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11416__A3 (.I(_01799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11417__B (.I(_00512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11418__A1 (.I(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11418__B (.I(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11418__C (.I(_00541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11419__A2 (.I(_00788_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11419__B (.I(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11420__A1 (.I(_02536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11421__A2 (.I(_01801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11421__A3 (.I(_03729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11422__A1 (.I(_04048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11423__A1 (.I(_02538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11425__A3 (.I(_04397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11426__I (.I(_05477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11427__A1 (.I(_04033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11428__A1 (.I(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11429__B (.I(_00840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11430__A1 (.I(_04240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11430__C (.I(_02173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11431__B (.I(_00773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11448__A3 (.I(_02246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11449__I (.I(_05491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11451__I (.I(_05491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11452__A1 (.I(\as2650.stack[9][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11452__A2 (.I(_05494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11455__I (.I(_05497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11456__A1 (.I(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11457__I (.I(_05491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11459__A1 (.I(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11461__A1 (.I(_02692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11463__A1 (.I(_02694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11466__I (.I(_05497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11467__A1 (.I(_02696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11468__A1 (.I(\as2650.stack[9][13] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11469__A1 (.I(_02700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11470__A1 (.I(\as2650.stack[9][14] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11471__A1 (.I(_02702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11473__I (.I(_05508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11474__A3 (.I(_02253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11477__A1 (.I(_01840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11478__A1 (.I(_03557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11478__B2 (.I(_05513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11479__A1 (.I(\as2650.stack[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11480__I (.I(_05491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11481__I (.I(_05497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11482__A2 (.I(_05515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11482__B (.I(_05516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11483__A1 (.I(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11484__A1 (.I(\as2650.stack[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11485__A1 (.I(_01870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11485__A2 (.I(_05515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11485__B (.I(_05516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11486__A1 (.I(_03569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11487__A1 (.I(\as2650.stack[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11488__A1 (.I(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11488__A2 (.I(_05515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11488__B (.I(_05516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11489__A1 (.I(_03572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11490__I (.I(_05497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11492__A1 (.I(\as2650.stack[9][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11492__A2 (.I(_05523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11493__A1 (.I(_01892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11493__A2 (.I(_05515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11493__B (.I(_05516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11495__A1 (.I(\as2650.stack[9][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11495__A2 (.I(_05523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11496__A2 (.I(_05494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11496__B (.I(_05508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11497__A1 (.I(_03580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11498__A1 (.I(\as2650.stack[9][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11498__A2 (.I(_05523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11499__A2 (.I(_05494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11499__B (.I(_05508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11501__A1 (.I(\as2650.stack[9][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11501__A2 (.I(_05523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11502__A2 (.I(_05494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11502__B (.I(_05508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11504__A1 (.I(_00947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11506__A1 (.I(_00946_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11506__C (.I(_00909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11507__I (.I(_05534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11509__A2 (.I(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11509__B2 (.I(_01141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11510__I (.I(_01401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11512__A2 (.I(_03397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11512__B2 (.I(_01233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11514__A2 (.I(_03429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11514__B2 (.I(_01305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11516__A2 (.I(_03458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11516__B2 (.I(_01375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11518__I (.I(_05534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11520__A2 (.I(_03477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11520__B2 (.I(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11522__A2 (.I(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11522__B2 (.I(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11524__A2 (.I(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11524__B2 (.I(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11526__A2 (.I(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11526__B2 (.I(_01718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11527__I (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11530__I0 (.I(_01225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11530__I1 (.I(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11531__A1 (.I(_00631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11531__C (.I(_00477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11532__A1 (.I(_00627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11533__B (.I(_00884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11533__C (.I(_00635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11535__A1 (.I(_00876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11535__A2 (.I(_01180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11535__A3 (.I(_03858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11535__A4 (.I(_00501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11536__A3 (.I(_05555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11538__I (.I(_05557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11539__I1 (.I(_05550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11540__A1 (.I(_05042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11541__I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11544__A1 (.I(_01851_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11546__I1 (.I(_05564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11547__A1 (.I(_05042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11548__I0 (.I(_00441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11548__I1 (.I(_01865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11549__I0 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11549__I1 (.I(_05566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11550__A1 (.I(_02570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11552__I0 (.I(_05252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11552__I1 (.I(_02097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11553__I (.I(_05557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11554__I0 (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11554__I1 (.I(_05569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11555__A1 (.I(_02570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11557__I0 (.I(_05341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11557__I1 (.I(_01421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11558__I0 (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11558__I1 (.I(_05573_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11559__A1 (.I(_02570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11561__I (.I(_00846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11562__A1 (.I(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11563__A1 (.I(_01900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11564__I0 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11564__I1 (.I(_05578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11565__A1 (.I(_05576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11567__I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11568__A1 (.I(_01911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11569__A1 (.I(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11571__A1 (.I(_05042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11572__I0 (.I(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11572__I1 (.I(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11573__I0 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11573__I1 (.I(_05585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11574__A1 (.I(_05576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11592__A1 (.I(_02850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11593__A1 (.I(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11594__A1 (.I(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11595__A1 (.I(_00877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11596__A1 (.I(_00838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11596__A2 (.I(_02750_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11596__A3 (.I(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11598__A1 (.I(_00965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11600__A1 (.I(_01368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11603__A1 (.I(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11605__A1 (.I(_01117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11605__A2 (.I(_00675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11605__A3 (.I(_02798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11605__A4 (.I(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11606__A2 (.I(_02565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11606__B1 (.I(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11608__A1 (.I(_04640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11608__A3 (.I(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11609__A1 (.I(_01063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11609__B (.I(_01065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11610__A1 (.I(_00919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11610__A2 (.I(_02565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11610__A3 (.I(_01063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11614__A2 (.I(_04460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11615__A1 (.I(_05615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11618__B (.I(_01157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11620__A1 (.I(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11621__A1 (.I(_01225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11622__A1 (.I(_02549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11622__A2 (.I(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11622__B (.I(_04461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11623__A1 (.I(_02896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11623__C (.I(_00963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11624__A1 (.I(_00628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11625__B (.I(_05408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11626__A2 (.I(_04585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11627__A1 (.I(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11627__C (.I(_05088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11628__A2 (.I(_01965_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11630__A1 (.I(_00839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11630__A2 (.I(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11631__A1 (.I(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11633__A1 (.I(_00583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11634__I (.I(_01787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11635__A1 (.I(_01324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11635__B (.I(_01929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11635__C (.I(_04885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11637__A1 (.I(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11638__A1 (.I(_04473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11638__A2 (.I(_00942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11638__B (.I(_04587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11639__I (.I(_02093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11640__A1 (.I(_02566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11640__B1 (.I(_05639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11640__B2 (.I(_05640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11640__C (.I(_00960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11641__A1 (.I(_05262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11642__A2 (.I(_05631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11642__B2 (.I(_04984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11643__A1 (.I(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11643__A2 (.I(_01003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11644__A1 (.I(_00969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11644__A2 (.I(_04587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11646__A1 (.I(_05477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11647__I1 (.I(_01785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11648__A1 (.I(_05576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11650__A2 (.I(_04559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11651__A1 (.I(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11651__A2 (.I(_01003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11651__A3 (.I(_05650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11651__B (.I(_05477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11652__A1 (.I(_02406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11652__A2 (.I(_02298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11654__A1 (.I(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11655__A1 (.I(_01271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11655__B (.I(_01929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11655__C (.I(_04885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11657__A1 (.I(_02860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11658__A1 (.I(_02003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11658__A2 (.I(_05639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11658__B2 (.I(_02566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11658__C (.I(_00960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11659__A1 (.I(_05245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11660__A1 (.I(_05631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11660__B2 (.I(_04984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11662__A1 (.I(_02406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11662__C (.I(_05088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11663__A1 (.I(_04501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11663__A2 (.I(_01003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11666__A1 (.I(_01981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11666__A2 (.I(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11667__A1 (.I(_02547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11667__A2 (.I(_01798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11668__A1 (.I(_01209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11668__A2 (.I(_00974_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11668__B1 (.I(_00975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11668__B2 (.I(_05665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11668__C (.I(_00919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11669__A1 (.I(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11669__A2 (.I(_04467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11670__A1 (.I(_05282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11670__A2 (.I(_05227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11670__A3 (.I(_05639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11670__B2 (.I(_02566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11671__A2 (.I(_00839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11671__B1 (.I(_00960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11672__A1 (.I(_05665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11672__B2 (.I(_03981_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11674__A1 (.I(_01822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11674__C (.I(_04757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11675__A1 (.I(_00537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11675__A2 (.I(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11675__B (.I(_05615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11676__A1 (.I(_02497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11676__A2 (.I(_02550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11676__B (.I(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11677__A1 (.I(_05341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11679__A1 (.I(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11679__A2 (.I(_04824_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11679__B1 (.I(_05676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11679__C (.I(_05673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11682__A1 (.I(_00553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11682__A2 (.I(_05679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11683__A1 (.I(_01895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11683__A2 (.I(_05673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11684__A1 (.I(_00996_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11685__A1 (.I(_04718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11685__A2 (.I(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11687__I (.I(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11688__A1 (.I(_01865_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11688__A2 (.I(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11688__B2 (.I(_04475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11690__A1 (.I(_05195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11690__A2 (.I(_04664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11691__A2 (.I(_03228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11692__A2 (.I(_03228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11692__C (.I(_00553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11693__A1 (.I(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11693__B2 (.I(_05689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11693__C (.I(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11694__A1 (.I(_00897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11694__A2 (.I(_00807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11694__A3 (.I(_04558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11697__A1 (.I(_04447_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11697__A2 (.I(_04801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11698__A1 (.I(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11698__A2 (.I(_00795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11698__C (.I(_00840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11699__A1 (.I(_05194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11699__A2 (.I(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11699__A3 (.I(_02850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11700__B (.I(_01230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11702__A1 (.I(_05576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11703__I (.I(_05698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11705__A1 (.I(_02097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11705__A2 (.I(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11706__A1 (.I(_00840_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11707__A1 (.I(_05195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11707__A2 (.I(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11708__A1 (.I(_01873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11708__C (.I(_04757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11710__A1 (.I(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11710__A2 (.I(_04501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11711__B (.I(_05408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11712__A1 (.I(_05195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11712__A2 (.I(_04612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11713__A1 (.I(_01846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11713__C (.I(_04757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11714__A1 (.I(_00795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11714__A2 (.I(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11715__A1 (.I(_03625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11715__A2 (.I(_04489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11715__B1 (.I(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11716__A1 (.I(_02343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11717__A1 (.I(_02343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11717__B (.I(_02923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11718__A1 (.I(_04702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11720__A1 (.I(_04489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11720__A2 (.I(_04003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11720__B (.I(_02343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11721__A1 (.I(_05725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11722__A1 (.I(_03622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11722__A2 (.I(_00538_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11723__A1 (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11723__B (.I(_00846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11789__CLK (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11790__CLK (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11850__CLK (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11888__CLK (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11952__CLK (.I(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11957__CLK (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__11999__CLK (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12012__CLK (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12018__D (.I(_00293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12039__D (.I(_00314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12044__CLK (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12047__CLK (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12054__D (.I(_00329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12055__D (.I(_00330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12057__D (.I(_00332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12076__D (.I(_00351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12077__D (.I(_00352_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12078__D (.I(_00353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12079__D (.I(_00354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12080__D (.I(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12081__D (.I(_00356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12089__CLK (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12090__CLK (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12091__CLK (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12114__CLK (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12121__CLK (.I(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12123__CLK (.I(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12129__CLK (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12130__CLK (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12134__D (.I(_00409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12138__CLK (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12141__D (.I(_00416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12223__I (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12224__I (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__12225__I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_wb_clk_i_I (.I(wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_0_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_1_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_2_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_3_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_4_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_5_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_6_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_7_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_0__f_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_10__f_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_11__f_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_12__f_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_13__f_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_14__f_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_15__f_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_1__f_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_2__f_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_3__f_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_4__f_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_5__f_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_6__f_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_7__f_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_8__f_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_4_9__f_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_0_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_100_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_102_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_103_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_104_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_105_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_106_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_107_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_109_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_10_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_111_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_112_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_113_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_114_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_115_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_116_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_117_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_118_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_119_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_11_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_120_wb_clk_i_I (.I(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_123_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_125_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_126_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_127_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_12_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_13_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_14_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_15_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_16_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_17_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_18_wb_clk_i_I (.I(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_19_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_1_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_20_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_21_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_22_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_23_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_24_wb_clk_i_I (.I(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_25_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_26_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_27_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_28_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_29_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_2_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_31_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_32_wb_clk_i_I (.I(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_33_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_34_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_35_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_36_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_37_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_38_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_39_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_3_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_40_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_41_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_42_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_43_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_44_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_46_wb_clk_i_I (.I(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_48_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_49_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_4_wb_clk_i_I (.I(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_50_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_52_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_53_wb_clk_i_I (.I(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_58_wb_clk_i_I (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_59_wb_clk_i_I (.I(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_5_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_60_wb_clk_i_I (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_61_wb_clk_i_I (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_63_wb_clk_i_I (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_64_wb_clk_i_I (.I(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_65_wb_clk_i_I (.I(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_66_wb_clk_i_I (.I(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_67_wb_clk_i_I (.I(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_68_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_69_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_6_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_70_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_71_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_72_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_73_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_74_wb_clk_i_I (.I(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_75_wb_clk_i_I (.I(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_76_wb_clk_i_I (.I(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_77_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_78_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_79_wb_clk_i_I (.I(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_7_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_81_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_82_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_83_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_84_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_85_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_86_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_87_wb_clk_i_I (.I(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_8_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_91_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_92_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_93_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_94_wb_clk_i_I (.I(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_95_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_96_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_97_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_98_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_99_wb_clk_i_I (.I(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_9_wb_clk_i_I (.I(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout100_I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout87_I (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout88_I (.I(net89));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout89_I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout91_I (.I(net67));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout92_I (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout93_I (.I(net63));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout94_I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout95_I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout96_I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout97_I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout98_I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout99_I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(io_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(io_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(io_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(io_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(io_in[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(io_in[33]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(io_in[34]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(io_in[35]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(io_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output15_I (.I(net88));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output21_I (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output22_I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output23_I (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output24_I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output25_I (.I(net25));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output26_I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output27_I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output28_I (.I(net28));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output29_I (.I(net29));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output30_I (.I(net30));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output31_I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output32_I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output33_I (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output34_I (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output35_I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output36_I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output37_I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output38_I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output39_I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output40_I (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output41_I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output42_I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output43_I (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output44_I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output45_I (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output46_I (.I(net46));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output47_I (.I(net47));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output48_I (.I(net90));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output49_I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output50_I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output51_I (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output52_I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output53_I (.I(net101));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output54_I (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output55_I (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output56_I (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output57_I (.I(net57));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output58_I (.I(net58));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output59_I (.I(net59));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output60_I (.I(net60));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output61_I (.I(net61));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output62_I (.I(net62));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output63_I (.I(net93));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output64_I (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output65_I (.I(net92));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output66_I (.I(net66));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output67_I (.I(net91));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output68_I (.I(net68));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output69_I (.I(net69));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output70_I (.I(net70));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output71_I (.I(net71));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output72_I (.I(net72));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output73_I (.I(net73));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output74_I (.I(net74));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output75_I (.I(net75));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output77_I (.I(net77));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output78_I (.I(net78));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output79_I (.I(net79));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire80_I (.I(_01304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire81_I (.I(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_wire82_I (.I(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_100_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_100_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_100_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_100_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_100_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_100_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_100_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_101_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_101_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_101_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_101_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_101_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_101_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_101_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_101_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_102_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_102_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_102_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_102_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_102_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_102_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_102_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_103_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_103_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_103_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_103_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_103_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_103_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_103_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_103_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_103_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_103_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_103_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_104_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_104_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_104_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_104_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_104_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_104_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_105_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_105_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_105_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_105_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_105_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_105_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_105_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_105_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_105_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_105_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_106_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_106_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_106_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_106_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_106_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_106_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_106_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_107_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_107_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_107_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_107_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_107_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_107_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_108_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_108_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_108_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_108_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_108_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_108_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_108_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_109_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_109_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_109_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_109_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_109_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_109_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_109_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_109_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_109_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_110_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_110_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_110_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_110_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_110_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_110_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_110_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_111_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_111_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_111_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_111_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_111_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_111_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_111_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_111_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_111_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_111_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_111_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_112_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_112_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_112_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_112_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_112_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_112_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_112_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_112_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_112_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_113_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_113_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_113_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_113_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_113_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_113_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_113_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_113_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_113_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_113_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_114_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_114_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_114_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_114_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_114_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_114_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_114_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_115_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_115_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_115_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_115_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_115_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_115_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_115_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_115_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_116_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_116_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_116_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_116_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_116_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_116_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_116_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_116_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_117_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_117_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_117_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_117_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_117_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_117_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_117_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_117_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_117_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_118_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_118_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_118_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_118_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_118_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_118_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_118_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_119_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_119_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_119_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_119_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_119_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_119_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_119_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_119_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_120_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_120_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_120_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_120_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_120_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_120_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_120_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_121_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_121_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_121_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_121_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_121_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_121_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_121_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_121_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_122_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_122_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_122_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_122_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_122_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_122_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_122_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_123_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_123_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_123_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_123_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_123_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_123_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_123_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_123_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_123_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_124_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_124_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_124_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_124_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_124_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_124_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_124_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_125_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_125_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_125_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_125_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_125_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_125_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_125_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_125_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_125_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_125_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_126_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_126_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_126_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_126_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_126_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_126_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_127_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_127_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_127_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_127_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_127_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_127_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_127_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_127_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_127_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_127_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_128_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_128_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_128_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_128_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_128_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_128_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_129_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_129_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_129_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_129_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_129_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_129_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_129_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_129_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_130_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_130_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_130_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_130_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_130_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_130_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_130_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_131_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_131_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_131_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_131_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_131_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_131_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_132_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_132_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_132_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_132_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_132_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_132_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_132_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_133_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_133_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_133_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_133_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_133_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_133_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_133_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_134_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_134_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_134_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_134_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_134_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_134_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_134_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_135_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_135_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_135_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_135_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_135_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_135_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_135_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_136_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_136_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_136_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_136_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_136_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_136_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_136_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_137_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_137_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_137_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_137_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_137_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_137_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_137_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_137_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_137_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_138_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_138_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_138_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_138_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_138_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_138_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_138_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_139_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_139_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_139_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_139_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_139_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_139_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_139_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_139_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_139_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_139_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_139_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_140_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_140_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_140_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_140_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_140_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_140_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_140_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_141_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_141_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_141_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_141_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_141_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_141_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_141_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_141_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_141_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_142_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_142_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_142_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_142_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_142_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_142_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_143_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_143_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_143_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_143_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_143_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_143_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_143_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_143_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_143_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_143_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_143_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_143_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_144_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_144_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_144_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_144_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_144_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_144_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_144_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_145_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_145_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_145_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_145_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_145_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_145_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_145_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_145_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_145_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_146_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_146_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_146_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_146_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_146_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_146_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_146_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_146_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_147_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_147_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_147_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_147_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_147_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_147_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_147_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_147_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_148_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_148_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_148_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_148_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_148_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_148_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_148_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_148_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_148_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_148_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_148_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_148_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_148_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_149_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_149_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_149_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_149_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_149_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_149_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_149_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_149_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_149_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_149_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_149_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_150_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_150_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_150_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_150_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_150_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_150_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_150_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_150_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_150_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_150_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_150_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_151_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_151_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_151_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_151_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_151_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_151_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_151_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_151_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_151_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_151_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_151_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_152_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_152_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_152_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_152_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_152_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_152_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_152_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_152_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_153_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_153_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_153_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_153_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_153_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_153_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_153_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_153_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_153_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_153_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_154_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_154_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_154_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_154_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_154_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_154_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_154_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_154_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_154_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_155_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_155_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_155_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_155_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_155_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_155_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_155_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_155_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_156_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_156_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_156_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_156_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_156_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_156_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_156_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_157_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_157_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_157_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_157_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_157_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_157_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_157_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_157_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_157_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_157_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_158_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_158_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_158_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_158_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_158_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_158_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_158_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_158_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_158_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_158_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_158_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_159_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_159_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_159_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_159_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_159_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_159_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_159_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_159_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_160_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_160_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_160_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_160_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_160_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_160_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_160_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_160_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_160_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_161_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_161_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_161_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_161_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_161_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_161_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_161_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_161_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_161_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_161_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_161_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_161_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_161_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_161_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_161_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_161_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_161_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_161_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_161_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_161_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_162_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_162_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_162_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_162_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_162_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_162_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_162_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_162_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_162_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_162_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_162_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_162_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_162_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_162_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_162_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_162_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_162_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_163_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_163_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_163_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_163_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_163_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_163_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_163_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_163_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_163_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_163_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_163_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_163_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_163_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_163_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_163_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_163_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_163_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_164_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_164_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_164_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_164_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_164_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_164_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_164_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_164_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_164_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_164_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_165_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_165_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_165_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_165_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_165_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_165_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_165_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_165_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_165_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_166_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_166_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_166_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_166_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_166_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_166_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_166_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_166_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_167_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_167_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_167_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_167_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_167_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_167_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_167_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_167_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_168_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_168_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_168_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_168_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_168_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_168_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_168_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_169_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_169_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_169_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_169_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_169_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_169_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_169_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_170_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_170_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_170_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_170_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_170_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_170_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_171_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_171_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_171_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_171_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_171_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_172_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_172_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_172_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_172_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_172_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_172_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_173_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_173_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_173_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_173_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_173_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_174_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_174_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_174_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_174_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_174_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_175_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_175_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_175_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_175_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_175_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_176_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_176_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_176_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_176_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_176_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_176_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_177_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_177_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_177_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_177_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_178_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_178_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_178_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_178_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_178_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_178_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_179_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_179_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_179_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_179_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_179_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_180_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_180_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_180_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_180_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_180_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_180_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_181_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_181_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_181_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_181_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_181_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_182_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_182_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_182_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_182_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_182_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_182_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_183_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_183_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_183_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_183_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_183_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_184_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_184_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_184_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_184_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_184_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_184_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_184_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_185_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_185_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_185_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_185_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_185_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_186_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_186_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_186_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_186_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_186_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_186_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_186_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_187_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_187_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_187_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_187_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_187_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_188_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_188_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_188_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_188_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_188_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_188_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_188_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_189_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_189_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_189_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_189_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_189_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_190_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_190_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_190_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_190_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_190_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_190_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_190_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_191_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_191_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_191_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_191_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_191_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_192_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_192_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_192_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_192_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_192_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_192_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_192_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_193_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_193_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_193_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_193_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_193_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_193_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_193_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_193_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_193_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_193_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_193_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_193_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_193_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_193_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_193_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_193_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_193_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_193_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_193_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_193_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_193_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_193_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_193_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_193_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_193_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_193_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_193_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_193_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_193_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_193_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_193_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_193_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_193_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_193_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_193_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_193_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_193_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_193_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_193_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_194_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_194_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_194_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_194_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_194_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_194_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_194_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_194_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_194_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_194_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_194_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_194_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_194_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_194_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_194_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_194_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_194_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_194_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_194_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_194_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_194_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_194_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_194_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_194_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_194_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_194_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_194_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_194_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_194_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_194_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_194_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_194_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_194_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_194_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_194_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_194_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_194_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_194_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_194_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_194_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_194_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_194_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_194_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_194_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_195_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_195_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_195_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_195_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_195_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_195_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_195_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_195_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_195_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_195_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_195_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_195_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_195_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_195_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_195_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_195_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_195_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_195_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_195_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_195_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_195_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_195_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_195_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_195_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_195_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_195_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_195_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_23_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_31_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_57_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_63_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_65_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_66_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_67_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_67_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_68_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_68_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_68_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_68_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_68_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_68_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_69_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_69_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_69_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_69_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_69_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_70_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_70_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_70_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_70_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_70_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_70_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_70_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_71_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_71_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_71_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_71_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_71_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_71_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_72_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_72_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_72_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_72_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_72_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_72_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_73_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_73_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_73_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_73_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_73_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_73_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_74_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_74_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_74_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_74_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_74_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_74_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_75_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_75_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_75_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_75_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_75_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_75_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_75_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_76_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_76_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_76_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_76_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_76_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_76_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_76_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_77_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_77_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_77_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_77_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_77_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_77_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_78_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_78_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_78_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_78_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_78_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_78_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_78_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_79_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_79_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_79_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_79_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_79_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_79_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_80_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_80_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_80_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_80_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_80_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_80_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_80_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_81_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_81_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_81_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_81_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_81_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_82_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_82_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_82_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_82_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_82_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_82_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_82_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_83_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_83_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_83_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_83_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_83_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_83_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_84_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_84_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_84_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_84_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_84_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_85_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_85_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_85_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_85_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_85_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_85_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_85_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_86_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_86_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_86_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_86_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_86_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_86_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_86_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_87_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_87_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_87_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_87_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_87_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_87_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_88_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_88_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_88_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_88_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_88_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_88_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_88_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_89_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_89_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_89_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_89_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_89_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_89_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_89_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_90_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_90_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_90_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_90_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_90_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_90_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_90_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_90_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_90_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_91_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_91_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_91_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_91_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_91_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_91_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_91_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_92_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_92_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_92_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_92_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_92_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_92_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_92_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_93_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_93_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_93_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_93_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_93_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_93_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_93_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_94_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_94_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_94_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_94_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_94_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_94_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_94_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_95_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_95_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_95_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_95_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_95_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_95_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_95_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_95_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_95_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_96_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_96_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_96_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_96_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_96_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_96_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_96_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_97_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_97_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_97_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_97_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_97_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_97_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_97_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_98_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_98_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_98_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_98_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_98_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_98_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_99_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_99_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_99_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_99_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_99_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_99_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_99_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_982 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_Left_296 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_100_Right_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_Left_297 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_101_Right_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_Left_298 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_102_Right_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_Left_299 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_103_Right_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_Left_300 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_104_Right_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_Left_301 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_105_Right_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_Left_302 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_106_Right_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_Left_303 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_107_Right_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_Left_304 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_108_Right_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_Left_305 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_109_Right_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_Left_306 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_110_Right_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_Left_307 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_111_Right_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_Left_308 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_112_Right_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_Left_309 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_113_Right_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_Left_310 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_114_Right_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_Left_311 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_115_Right_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_Left_312 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_116_Right_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_Left_313 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_117_Right_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_Left_314 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_118_Right_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_Left_315 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_119_Right_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_Left_316 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_120_Right_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_Left_317 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_121_Right_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_Left_318 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_122_Right_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_Left_319 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_123_Right_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_Left_320 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_124_Right_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_Left_321 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_125_Right_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_Left_322 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_126_Right_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_Left_323 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_127_Right_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_Left_324 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_128_Right_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_Left_325 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_129_Right_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_Left_326 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_130_Right_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_Left_327 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_131_Right_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_Left_328 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_132_Right_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_Left_329 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_133_Right_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_Left_330 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_134_Right_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_Left_331 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_135_Right_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_Left_332 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_136_Right_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_Left_333 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_137_Right_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_Left_334 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_138_Right_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_Left_335 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_139_Right_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_Left_336 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_140_Right_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_Left_337 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_141_Right_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_Left_338 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_142_Right_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_Left_339 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_143_Right_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_Left_340 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_144_Right_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_Left_341 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_145_Right_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_Left_342 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_146_Right_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_Left_343 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_147_Right_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_Left_344 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_148_Right_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_Left_345 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_149_Right_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_Left_346 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_150_Right_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_Left_347 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_151_Right_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_Left_348 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_152_Right_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_Left_349 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_153_Right_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_Left_350 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_154_Right_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_Left_351 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_155_Right_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_Left_352 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_156_Right_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_Left_353 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_157_Right_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_Left_354 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_158_Right_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_Left_355 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_159_Right_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_Left_356 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_160_Right_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_Left_357 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_161_Right_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_Left_358 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_162_Right_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_Left_359 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_163_Right_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_Left_360 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_164_Right_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_Left_361 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_165_Right_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_Left_362 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_166_Right_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_Left_363 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_167_Right_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_Left_364 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_168_Right_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_Left_365 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_169_Right_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_Left_366 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_170_Right_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_Left_367 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_171_Right_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_Left_368 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_172_Right_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_Left_369 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_173_Right_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_Left_370 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_174_Right_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_Left_371 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_175_Right_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_Left_372 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_176_Right_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_Left_373 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_177_Right_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_Left_374 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_178_Right_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_Left_375 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_179_Right_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_Left_376 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_180_Right_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_Left_377 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_181_Right_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_Left_378 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_182_Right_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_183_Left_379 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_183_Right_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_184_Left_380 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_184_Right_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_185_Left_381 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_185_Right_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_186_Left_382 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_186_Right_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_187_Left_383 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_187_Right_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_188_Left_384 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_188_Right_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_189_Left_385 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_189_Right_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_190_Left_386 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_190_Right_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_191_Left_387 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_191_Right_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_192_Left_388 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_192_Right_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_193_Left_389 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_193_Right_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_194_Left_390 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_194_Right_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_195_Left_391 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_195_Right_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Left_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Left_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Left_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Left_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Left_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Left_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Left_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Left_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Left_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Left_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Left_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Left_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Left_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Left_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Left_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Left_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Left_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Left_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Right_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Left_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Right_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Left_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Right_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Left_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Right_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Left_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Right_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Left_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Right_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Left_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_68_Right_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Left_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_69_Right_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Left_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_70_Right_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Left_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_71_Right_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Left_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_72_Right_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Left_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_73_Right_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Left_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_74_Right_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Left_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_75_Right_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Left_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_76_Right_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Left_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_77_Right_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Left_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_78_Right_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Left_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_79_Right_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Left_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_80_Right_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_Left_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_81_Right_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_Left_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_82_Right_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Left_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_83_Right_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Left_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_84_Right_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Left_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_85_Right_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Left_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_86_Right_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_Left_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_87_Right_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_Left_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_88_Right_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_Left_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_89_Right_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_Left_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_90_Right_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_Left_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_91_Right_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_Left_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_92_Right_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_Left_289 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_93_Right_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_Left_290 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_94_Right_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_Left_291 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_95_Right_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_Left_292 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_96_Right_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_Left_293 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_97_Right_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_Left_294 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_98_Right_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_Left_295 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_99_Right_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_100_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_101_3224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_102_3252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_103_3279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_104_3307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_105_3334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_106_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_107_3389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_108_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_109_3444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_110_3472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_111_3499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_112_3527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_113_3554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_114_3582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_115_3609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_116_3637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_117_3664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_118_3692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_119_3719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_120_3747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_121_3774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_122_3802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_123_3829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_124_3857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_125_3884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_126_3912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_127_3939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_128_3967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_129_3994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_3999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_130_4022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_131_4049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_132_4077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_133_4104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_134_4132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_135_4159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_136_4187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_137_4214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_138_4242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_139_4269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_140_4297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_141_4324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_142_4352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_143_4379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_144_4407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_145_4434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_146_4462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_147_4489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_148_4517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_149_4544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_150_4572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_151_4599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_152_4627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_153_4654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_154_4682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_155_4709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_156_4737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_157_4764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_158_4792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_159_4819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_160_4847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_161_4874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_162_4902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_163_4929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_164_4957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_165_4984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_4999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_5000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_5001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_5002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_5003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_5004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_5005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_5006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_5007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_5008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_5009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_5010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_5011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_166_5012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_167_5039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_168_5067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_169_5094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_170_5122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_171_5149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_172_5177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_173_5204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_174_5232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_175_5259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_176_5287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_177_5314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_178_5342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_179_5369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_180_5397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_181_5424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_182_5452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_183_5479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_184_5507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_185_5534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_186_5562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_187_5589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_188_5617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_189_5644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_190_5672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_191_5699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_192_5727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_193_5754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_194_5782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_195_5838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_68_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_69_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_70_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_71_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_72_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_73_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_74_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_75_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_76_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_77_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_78_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_79_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_80_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_81_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_82_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_83_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_84_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_85_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_86_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_87_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_88_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_89_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_90_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_91_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_92_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_93_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_94_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_95_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_96_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_97_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_98_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_99_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_694 ();
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05862_ (.I(net5),
    .Z(_05716_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05863_ (.I(_05716_),
    .Z(_05717_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05864_ (.I(_05717_),
    .Z(_05718_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05865_ (.I(_05718_),
    .Z(_05719_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05866_ (.I(\as2650.ins_reg[4] ),
    .ZN(_05720_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05867_ (.I(_05720_),
    .Z(_05721_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05868_ (.I(net54),
    .Z(_05722_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05869_ (.I(\as2650.ins_reg[1] ),
    .Z(_05723_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05870_ (.I(_05723_),
    .ZN(_05724_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05871_ (.I(_05724_),
    .Z(_05725_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05872_ (.A1(_05722_),
    .A2(_05725_),
    .ZN(_05726_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _05873_ (.I(net54),
    .ZN(_05727_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05874_ (.I(_05723_),
    .Z(_05728_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05875_ (.A1(_05727_),
    .A2(_05728_),
    .ZN(_05729_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05876_ (.I(\as2650.ins_reg[0] ),
    .Z(_05730_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05877_ (.I(_05730_),
    .Z(_05731_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05878_ (.I(_05731_),
    .Z(_05732_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _05879_ (.I(_05732_),
    .ZN(_05733_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05880_ (.A1(net101),
    .A2(_05733_),
    .ZN(_05734_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05881_ (.I(net101),
    .ZN(_05735_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05882_ (.I(_05732_),
    .Z(_05736_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05883_ (.A1(_05735_),
    .A2(_05736_),
    .ZN(_05737_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _05884_ (.A1(_05726_),
    .A2(_05729_),
    .A3(_05734_),
    .A4(_05737_),
    .ZN(_05738_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05885_ (.I(\as2650.alu_op[2] ),
    .Z(_05739_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05886_ (.I(_05739_),
    .Z(_05740_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05887_ (.I(\as2650.alu_op[1] ),
    .Z(_05741_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _05888_ (.I(_05741_),
    .ZN(_05742_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05889_ (.A1(_05740_),
    .A2(_05742_),
    .ZN(_05743_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05890_ (.I(_05743_),
    .Z(_05744_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05891_ (.A1(_05728_),
    .A2(_05736_),
    .ZN(_05745_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05892_ (.A1(_05745_),
    .A2(_05738_),
    .ZN(_05746_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05893_ (.I(\as2650.ins_reg[4] ),
    .Z(_05747_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05894_ (.A1(_05739_),
    .A2(_05741_),
    .ZN(_05748_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _05895_ (.A1(_05747_),
    .A2(_05748_),
    .ZN(_05749_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _05896_ (.A1(_05721_),
    .A2(_05738_),
    .A3(_05744_),
    .B1(_05746_),
    .B2(_05749_),
    .ZN(_05750_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05897_ (.I(net84),
    .ZN(_05751_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05898_ (.I(\as2650.ins_reg[4] ),
    .Z(_05752_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05899_ (.I(_05752_),
    .Z(_05753_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _05900_ (.I(_05753_),
    .Z(_05754_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05901_ (.I(_05741_),
    .Z(_05755_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _05902_ (.I(_05755_),
    .Z(_05756_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05903_ (.I(\as2650.r0[7] ),
    .Z(_05757_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05904_ (.I(_05757_),
    .Z(_05758_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _05905_ (.A1(_05723_),
    .A2(_05730_),
    .ZN(_05759_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05906_ (.I(_05759_),
    .Z(_05760_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05907_ (.I(_05760_),
    .Z(_05761_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05908_ (.I(_05761_),
    .Z(_05762_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _05909_ (.A1(_05728_),
    .A2(_05733_),
    .ZN(_05763_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05910_ (.I(net51),
    .Z(_05764_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05911_ (.I0(\as2650.r123[0][7] ),
    .I1(\as2650.r123_2[0][7] ),
    .S(_05764_),
    .Z(_05765_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05912_ (.I(_05765_),
    .Z(_05766_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05913_ (.I(_05766_),
    .Z(_05767_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _05914_ (.A1(_05758_),
    .A2(_05762_),
    .B1(_05763_),
    .B2(_05767_),
    .ZN(_05768_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05915_ (.A1(\as2650.ins_reg[1] ),
    .A2(_05730_),
    .Z(_05769_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05916_ (.I(_05769_),
    .Z(_05770_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05917_ (.I(_05770_),
    .Z(_05771_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05918_ (.I(_05771_),
    .Z(_05772_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _05919_ (.I(_05772_),
    .Z(_05773_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05920_ (.I(net51),
    .Z(_05774_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05921_ (.I(_05774_),
    .Z(_05775_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05922_ (.I(_05775_),
    .Z(_05776_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05923_ (.I(_05776_),
    .Z(_05777_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _05924_ (.I0(\as2650.r123[2][7] ),
    .I1(\as2650.r123_2[2][7] ),
    .S(_05777_),
    .Z(_05778_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05925_ (.A1(_05773_),
    .A2(_05778_),
    .ZN(_05779_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05926_ (.I(_05777_),
    .Z(_05780_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _05927_ (.I(_05780_),
    .ZN(_05781_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05928_ (.A1(_05724_),
    .A2(_05736_),
    .ZN(_05782_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05929_ (.A1(_05780_),
    .A2(\as2650.r123[1][7] ),
    .Z(_05783_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _05930_ (.A1(_05781_),
    .A2(\as2650.r123_2[1][7] ),
    .B(_05782_),
    .C(_05783_),
    .ZN(_05784_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _05931_ (.A1(_05768_),
    .A2(_05779_),
    .A3(_05784_),
    .Z(_05785_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05932_ (.I(\as2650.r0[5] ),
    .Z(_05786_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05933_ (.I(_05786_),
    .Z(_05787_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05934_ (.A1(_05787_),
    .A2(_05761_),
    .ZN(_05788_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05935_ (.I0(\as2650.r123[2][5] ),
    .I1(\as2650.r123_2[2][5] ),
    .S(_05776_),
    .Z(_05789_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _05936_ (.I0(\as2650.r123[1][5] ),
    .I1(\as2650.r123[0][5] ),
    .I2(\as2650.r123_2[1][5] ),
    .I3(\as2650.r123_2[0][5] ),
    .S0(_05731_),
    .S1(_05776_),
    .Z(_05790_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _05937_ (.A1(\as2650.ins_reg[1] ),
    .A2(\as2650.ins_reg[0] ),
    .Z(_05791_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05938_ (.I(_05791_),
    .Z(_05792_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05939_ (.I(_05792_),
    .Z(_05793_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _05940_ (.A1(_05771_),
    .A2(_05789_),
    .B1(_05790_),
    .B2(_05793_),
    .ZN(_05794_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05941_ (.A1(_05788_),
    .A2(_05794_),
    .Z(_05795_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05942_ (.I(\as2650.r0[4] ),
    .Z(_05796_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05943_ (.I(_05796_),
    .Z(_05797_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05944_ (.A1(_05797_),
    .A2(_05760_),
    .ZN(_05798_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05945_ (.I(_05774_),
    .Z(_05799_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05946_ (.I(_05799_),
    .Z(_05800_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _05947_ (.I0(\as2650.r123[2][4] ),
    .I1(\as2650.r123_2[2][4] ),
    .S(_05800_),
    .Z(_05801_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _05948_ (.I0(\as2650.r123[1][4] ),
    .I1(\as2650.r123[0][4] ),
    .I2(\as2650.r123_2[1][4] ),
    .I3(\as2650.r123_2[0][4] ),
    .S0(_05731_),
    .S1(_05800_),
    .Z(_05802_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _05949_ (.A1(_05770_),
    .A2(_05801_),
    .B1(_05802_),
    .B2(_05792_),
    .ZN(_05803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05950_ (.A1(_05798_),
    .A2(_05803_),
    .ZN(_05804_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05951_ (.I(_05804_),
    .Z(_05805_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05952_ (.I(\as2650.r0[3] ),
    .Z(_05806_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05953_ (.I(_05806_),
    .Z(_05807_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05954_ (.I(_05807_),
    .Z(_05808_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05955_ (.I(_05808_),
    .Z(_05809_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05956_ (.A1(_05809_),
    .A2(_05761_),
    .ZN(_05810_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _05957_ (.I0(\as2650.r123[2][3] ),
    .I1(\as2650.r123_2[2][3] ),
    .S(_05776_),
    .Z(_05811_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _05958_ (.I0(\as2650.r123[1][3] ),
    .I1(\as2650.r123[0][3] ),
    .I2(\as2650.r123_2[1][3] ),
    .I3(\as2650.r123_2[0][3] ),
    .S0(_05731_),
    .S1(_05800_),
    .Z(_05812_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _05959_ (.A1(_05771_),
    .A2(_05811_),
    .B1(_05812_),
    .B2(_05793_),
    .ZN(_05813_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05960_ (.A1(_05810_),
    .A2(_05813_),
    .ZN(_05814_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05961_ (.I(\as2650.r0[2] ),
    .Z(_05815_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _05962_ (.I(_05815_),
    .Z(_05816_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05963_ (.I(_05816_),
    .Z(_05817_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _05964_ (.I0(\as2650.r123[1][2] ),
    .I1(\as2650.r123[0][2] ),
    .I2(\as2650.r123_2[1][2] ),
    .I3(\as2650.r123_2[0][2] ),
    .S0(_05730_),
    .S1(_05775_),
    .Z(_05818_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _05965_ (.I0(\as2650.r123[2][2] ),
    .I1(\as2650.r123_2[2][2] ),
    .S(_05800_),
    .Z(_05819_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _05966_ (.A1(_05817_),
    .A2(_05760_),
    .B1(_05792_),
    .B2(_05818_),
    .C1(_05819_),
    .C2(_05770_),
    .ZN(_05820_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05967_ (.I(_05820_),
    .Z(_05821_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05968_ (.I(_05821_),
    .Z(_05822_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _05969_ (.I(\as2650.r0[1] ),
    .Z(_05823_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05970_ (.I(_05823_),
    .Z(_05824_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _05971_ (.I0(\as2650.r123[1][1] ),
    .I1(\as2650.r123[0][1] ),
    .I2(\as2650.r123_2[1][1] ),
    .I3(\as2650.r123_2[0][1] ),
    .S0(\as2650.ins_reg[0] ),
    .S1(_05775_),
    .Z(_05825_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _05972_ (.I0(\as2650.r123[2][1] ),
    .I1(\as2650.r123_2[2][1] ),
    .S(_05775_),
    .Z(_05826_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _05973_ (.A1(_05824_),
    .A2(_05759_),
    .B1(_05792_),
    .B2(_05825_),
    .C1(_05826_),
    .C2(_05770_),
    .ZN(_05827_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05974_ (.I(_05827_),
    .Z(_05828_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _05975_ (.A1(\as2650.ins_reg[4] ),
    .A2(\as2650.alu_op[2] ),
    .A3(\as2650.alu_op[1] ),
    .ZN(_05829_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05976_ (.I(\as2650.r0[0] ),
    .Z(_05830_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_4 _05977_ (.I0(\as2650.r123[1][0] ),
    .I1(\as2650.r123[0][0] ),
    .I2(\as2650.r123_2[1][0] ),
    .I3(\as2650.r123_2[0][0] ),
    .S0(\as2650.ins_reg[0] ),
    .S1(_05799_),
    .Z(_05831_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _05978_ (.I0(\as2650.r123[2][0] ),
    .I1(\as2650.r123_2[2][0] ),
    .S(_05799_),
    .Z(_05832_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _05979_ (.A1(_05830_),
    .A2(_05759_),
    .B1(_05791_),
    .B2(_05831_),
    .C1(_05832_),
    .C2(_05769_),
    .ZN(_05833_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05980_ (.I(_05833_),
    .Z(_05834_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _05981_ (.A1(\as2650.alu_op[0] ),
    .A2(_05829_),
    .A3(_05834_),
    .Z(_05835_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _05982_ (.A1(_05822_),
    .A2(_05828_),
    .A3(_05835_),
    .ZN(_05836_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _05983_ (.A1(_05805_),
    .A2(_05814_),
    .A3(_05836_),
    .ZN(_05837_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05984_ (.A1(_05795_),
    .A2(_05837_),
    .Z(_05838_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _05985_ (.A1(_05788_),
    .A2(_05794_),
    .ZN(_05839_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _05986_ (.I(_05839_),
    .Z(_05840_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05987_ (.I(_05833_),
    .Z(_05841_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05988_ (.I(\as2650.alu_op[0] ),
    .Z(_05842_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _05989_ (.I(_05842_),
    .ZN(_05843_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05990_ (.I(_05829_),
    .Z(_05844_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _05991_ (.A1(_05843_),
    .A2(_05844_),
    .ZN(_05845_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _05992_ (.A1(_05841_),
    .A2(_05845_),
    .ZN(_05846_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _05993_ (.A1(_05798_),
    .A2(_05803_),
    .Z(_05847_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05994_ (.I(_05847_),
    .Z(_05848_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _05995_ (.A1(_05809_),
    .A2(_05760_),
    .B1(_05793_),
    .B2(_05812_),
    .C1(_05811_),
    .C2(_05771_),
    .ZN(_05849_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _05996_ (.I(_05849_),
    .Z(_05850_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _05997_ (.A1(_05848_),
    .A2(_05850_),
    .A3(_05822_),
    .A4(_05828_),
    .ZN(_05851_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05998_ (.A1(_05846_),
    .A2(_05851_),
    .Z(_05852_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _05999_ (.A1(_05840_),
    .A2(_05852_),
    .Z(_05853_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06000_ (.I(\as2650.r0[6] ),
    .Z(_05854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06001_ (.I(_05854_),
    .Z(_05855_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06002_ (.A1(_05855_),
    .A2(_05761_),
    .ZN(_05856_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_4 _06003_ (.I0(\as2650.r123[2][6] ),
    .I1(\as2650.r123_2[2][6] ),
    .S(_05777_),
    .Z(_05857_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_2 _06004_ (.I0(\as2650.r123[1][6] ),
    .I1(\as2650.r123[0][6] ),
    .I2(\as2650.r123_2[1][6] ),
    .I3(\as2650.r123_2[0][6] ),
    .S0(_05732_),
    .S1(_05777_),
    .Z(_05858_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06005_ (.I(_05793_),
    .Z(_05859_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _06006_ (.A1(_05772_),
    .A2(_05857_),
    .B1(_05858_),
    .B2(_05859_),
    .ZN(_05860_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06007_ (.A1(_05856_),
    .A2(_05860_),
    .Z(_05861_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06008_ (.I0(_05838_),
    .I1(_05853_),
    .S(_05861_),
    .Z(_00420_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06009_ (.A1(_05785_),
    .A2(_00420_),
    .Z(_00421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06010_ (.A1(_05856_),
    .A2(_05860_),
    .ZN(_00422_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06011_ (.A1(_05838_),
    .A2(_05853_),
    .ZN(_00423_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06012_ (.A1(_00422_),
    .A2(_00423_),
    .Z(_00424_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06013_ (.I(_05840_),
    .Z(_00425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06014_ (.A1(_00425_),
    .A2(_05852_),
    .ZN(_00426_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06015_ (.A1(_05837_),
    .A2(_05853_),
    .A3(_00426_),
    .ZN(_00427_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _06016_ (.A1(_05838_),
    .A2(_00427_),
    .Z(_00428_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06017_ (.I(_05848_),
    .Z(_00429_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06018_ (.I(_05821_),
    .Z(_00430_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06019_ (.I(_05828_),
    .Z(_00431_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06020_ (.A1(_00430_),
    .A2(_00431_),
    .ZN(_00432_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06021_ (.A1(_05814_),
    .A2(_05846_),
    .A3(_00432_),
    .ZN(_00433_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06022_ (.I(_05814_),
    .Z(_00434_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06023_ (.A1(_00434_),
    .A2(_05836_),
    .ZN(_00435_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _06024_ (.A1(_00429_),
    .A2(_00433_),
    .B(_05852_),
    .C(_00435_),
    .ZN(_00436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06025_ (.A1(_05837_),
    .A2(_00436_),
    .ZN(_00437_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06026_ (.I(_05817_),
    .Z(_00438_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06027_ (.A1(_00438_),
    .A2(_05762_),
    .ZN(_00439_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _06028_ (.A1(_05772_),
    .A2(_05819_),
    .B1(_05818_),
    .B2(_05859_),
    .ZN(_00440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06029_ (.A1(_00439_),
    .A2(_00440_),
    .ZN(_00441_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06030_ (.I(_00431_),
    .Z(_00442_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06031_ (.I(_05834_),
    .Z(_00443_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06032_ (.I(_00443_),
    .Z(_00444_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06033_ (.I(_00444_),
    .Z(_00445_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06034_ (.A1(_00442_),
    .A2(_00445_),
    .A3(_05845_),
    .ZN(_00446_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06035_ (.A1(_05846_),
    .A2(_00432_),
    .ZN(_00447_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06036_ (.A1(_00442_),
    .A2(_05835_),
    .ZN(_00448_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06037_ (.A1(_00441_),
    .A2(_00446_),
    .B(_00447_),
    .C(_00448_),
    .ZN(_00449_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _06038_ (.A1(_05836_),
    .A2(_00449_),
    .Z(_00450_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06039_ (.A1(_05850_),
    .A2(_00447_),
    .ZN(_00451_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _06040_ (.A1(_05836_),
    .A2(_00433_),
    .A3(_00451_),
    .B(_00435_),
    .ZN(_00452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06041_ (.A1(_05835_),
    .A2(_05846_),
    .ZN(_00453_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06042_ (.A1(_00442_),
    .A2(_00453_),
    .Z(_00454_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _06043_ (.A1(_05844_),
    .A2(_00445_),
    .ZN(_00455_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _06044_ (.A1(_00450_),
    .A2(_00452_),
    .A3(_00454_),
    .A4(_00455_),
    .Z(_00456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06045_ (.A1(_00437_),
    .A2(_00456_),
    .ZN(_00457_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06046_ (.A1(_00421_),
    .A2(_00424_),
    .A3(_00428_),
    .A4(_00457_),
    .ZN(_00458_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06047_ (.A1(_05754_),
    .A2(_05756_),
    .A3(_00458_),
    .ZN(_00459_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06048_ (.A1(_05751_),
    .A2(_00459_),
    .ZN(_00460_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06049_ (.I(_00460_),
    .Z(_00461_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06050_ (.I(_00461_),
    .Z(_00462_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06051_ (.I(\as2650.ins_reg[3] ),
    .Z(_00463_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06052_ (.I(_00463_),
    .Z(_00464_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06053_ (.A1(_00464_),
    .A2(_05747_),
    .ZN(_00465_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06054_ (.I(_00465_),
    .Z(_00466_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06055_ (.I(_00466_),
    .Z(_00467_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06056_ (.I(_05739_),
    .ZN(_00468_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06057_ (.A1(_00468_),
    .A2(_05755_),
    .ZN(_00469_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _06058_ (.I(_00463_),
    .ZN(_00470_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06059_ (.A1(_00470_),
    .A2(_05720_),
    .ZN(_00471_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06060_ (.A1(_05773_),
    .A2(_00469_),
    .A3(_00471_),
    .ZN(_00472_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06061_ (.I(_00472_),
    .Z(_00473_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06062_ (.A1(_05723_),
    .A2(_05732_),
    .Z(_00474_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06063_ (.I(_00474_),
    .Z(_00475_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06064_ (.I(_05843_),
    .Z(_00476_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06065_ (.A1(_00476_),
    .A2(_05739_),
    .A3(_05741_),
    .ZN(_00477_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06066_ (.A1(_05752_),
    .A2(_00477_),
    .ZN(_00478_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06067_ (.I(\as2650.ins_reg[2] ),
    .Z(_00479_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06068_ (.I(_00479_),
    .ZN(_00480_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06069_ (.I(_00480_),
    .Z(_00481_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06070_ (.A1(_00481_),
    .A2(_00463_),
    .ZN(_00482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06071_ (.A1(_00478_),
    .A2(_00482_),
    .ZN(_00483_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06072_ (.A1(_00475_),
    .A2(_00483_),
    .ZN(_00484_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06073_ (.I(\as2650.prefixed ),
    .ZN(_00485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06074_ (.I(_00485_),
    .Z(_00486_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06075_ (.A1(net72),
    .A2(\as2650.cycle[0] ),
    .ZN(_00487_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06076_ (.I(_00487_),
    .Z(_00488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06077_ (.A1(_00486_),
    .A2(_00488_),
    .ZN(_00489_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06078_ (.A1(_00484_),
    .A2(_00489_),
    .ZN(_00490_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06079_ (.I(_00490_),
    .Z(_00491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06080_ (.A1(_00473_),
    .A2(_00491_),
    .ZN(_00492_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _06081_ (.A1(_05719_),
    .A2(_00462_),
    .A3(_00467_),
    .A4(_00492_),
    .ZN(_00493_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06082_ (.I(_05762_),
    .Z(_00494_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06083_ (.A1(_00494_),
    .A2(_00478_),
    .A3(_00482_),
    .ZN(_00495_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06084_ (.A1(_00495_),
    .A2(_00488_),
    .ZN(_00496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06085_ (.A1(_00486_),
    .A2(_00470_),
    .ZN(_00497_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06086_ (.A1(_00496_),
    .A2(_00497_),
    .ZN(_00498_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06087_ (.I(_05716_),
    .Z(_00499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06088_ (.A1(_05842_),
    .A2(_05752_),
    .ZN(_00500_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06089_ (.A1(_00479_),
    .A2(_00500_),
    .ZN(_00501_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06090_ (.A1(_05740_),
    .A2(_00501_),
    .ZN(_00502_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06091_ (.I(_00502_),
    .Z(_00503_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06092_ (.A1(_00499_),
    .A2(_00503_),
    .ZN(_00504_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06093_ (.A1(_00498_),
    .A2(_00504_),
    .Z(_00505_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06094_ (.I(_05717_),
    .Z(_00506_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06095_ (.I(_00506_),
    .Z(_00507_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06096_ (.I(_00479_),
    .Z(_00508_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06097_ (.I(_00508_),
    .Z(_00509_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06098_ (.A1(_05745_),
    .A2(_05743_),
    .A3(_00465_),
    .ZN(_00510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06099_ (.A1(_00509_),
    .A2(_00510_),
    .ZN(_00511_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06100_ (.I(_00511_),
    .Z(_00512_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06101_ (.I(_00512_),
    .Z(_00513_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06102_ (.I(_00513_),
    .Z(_00514_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06103_ (.I(_00488_),
    .Z(_00515_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06104_ (.A1(\as2650.prefixed ),
    .A2(_00470_),
    .A3(_05720_),
    .ZN(_00516_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06105_ (.A1(_00515_),
    .A2(_00516_),
    .ZN(_00517_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06106_ (.I(_00517_),
    .Z(_00518_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06107_ (.I(net5),
    .ZN(_00519_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06108_ (.A1(_00519_),
    .A2(_00487_),
    .ZN(_00520_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06109_ (.I(_05747_),
    .Z(_00521_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06110_ (.A1(\as2650.prefixed ),
    .A2(_00464_),
    .ZN(_00522_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06111_ (.A1(_00521_),
    .A2(_00522_),
    .ZN(_00523_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06112_ (.A1(_00520_),
    .A2(_00523_),
    .ZN(_00524_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06113_ (.I(_05740_),
    .Z(_00525_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06114_ (.I(_00481_),
    .Z(_00526_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06115_ (.I(_05842_),
    .Z(_00527_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06116_ (.A1(_00526_),
    .A2(_00527_),
    .A3(_00521_),
    .ZN(_00528_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06117_ (.A1(_00525_),
    .A2(_00528_),
    .ZN(_00529_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06118_ (.A1(_00524_),
    .A2(_00529_),
    .ZN(_00530_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06119_ (.A1(_00507_),
    .A2(_00514_),
    .A3(_00518_),
    .B(_00530_),
    .ZN(_00531_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06120_ (.I(\as2650.cycle[6] ),
    .Z(_00532_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06121_ (.I(_00532_),
    .Z(_00533_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06122_ (.I(_00533_),
    .Z(_00534_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06123_ (.I(_00534_),
    .Z(_00535_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06124_ (.I(_00535_),
    .Z(_00536_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06125_ (.I(_00536_),
    .Z(_00537_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06126_ (.I(_00537_),
    .Z(_00538_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06127_ (.A1(_00493_),
    .A2(_00505_),
    .A3(_00531_),
    .B(_00538_),
    .ZN(_00539_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06128_ (.A1(_00508_),
    .A2(_00472_),
    .ZN(_00540_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06129_ (.I(_00540_),
    .Z(_00541_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06130_ (.I(_00541_),
    .Z(_00542_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06131_ (.I(_00542_),
    .Z(_00543_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06132_ (.I(_00516_),
    .Z(_00544_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06133_ (.A1(_00515_),
    .A2(_00544_),
    .Z(_00545_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06134_ (.I(_00545_),
    .Z(_00546_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06135_ (.I(_00546_),
    .Z(_00547_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06136_ (.A1(_00543_),
    .A2(_00547_),
    .ZN(_00548_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06137_ (.I(\as2650.prefixed ),
    .Z(_00549_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06138_ (.A1(_00549_),
    .A2(_05753_),
    .ZN(_00550_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06139_ (.I(_00550_),
    .Z(_00551_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06140_ (.I(_00551_),
    .Z(_00552_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06141_ (.I(_00552_),
    .Z(_00553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06142_ (.A1(_00476_),
    .A2(_05752_),
    .ZN(_00554_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06143_ (.A1(_05743_),
    .A2(_00554_),
    .ZN(_00555_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06144_ (.A1(_00479_),
    .A2(_00463_),
    .ZN(_00556_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06145_ (.I(_00556_),
    .Z(_00557_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06146_ (.I(_00557_),
    .Z(_00558_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06147_ (.I(_00558_),
    .Z(_00559_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06148_ (.I(_00559_),
    .Z(_00560_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06149_ (.A1(_00494_),
    .A2(_00555_),
    .A3(_00560_),
    .ZN(_00561_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06150_ (.A1(_00485_),
    .A2(_05753_),
    .ZN(_00562_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06151_ (.A1(_00481_),
    .A2(_05749_),
    .ZN(_00563_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06152_ (.A1(_00464_),
    .A2(_00562_),
    .A3(_00563_),
    .ZN(_00564_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06153_ (.A1(_00515_),
    .A2(_00561_),
    .A3(_00564_),
    .ZN(_00565_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06154_ (.I(_00554_),
    .Z(_00566_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06155_ (.A1(_00468_),
    .A2(_05755_),
    .ZN(_00567_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06156_ (.A1(_00508_),
    .A2(_00566_),
    .A3(_00567_),
    .ZN(_00568_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06157_ (.A1(_00508_),
    .A2(_00527_),
    .A3(_05844_),
    .ZN(_00569_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06158_ (.A1(_00568_),
    .A2(_00569_),
    .ZN(_00570_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06159_ (.A1(_00528_),
    .A2(_00570_),
    .ZN(_00571_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06160_ (.A1(_00565_),
    .A2(_00571_),
    .ZN(_00572_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06161_ (.A1(net72),
    .A2(\as2650.cycle[0] ),
    .Z(_00573_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06162_ (.I(_00573_),
    .Z(_00574_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06163_ (.A1(_00484_),
    .A2(_00574_),
    .ZN(_00575_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06164_ (.I(_00575_),
    .Z(_00576_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _06165_ (.A1(_00553_),
    .A2(_00572_),
    .B(_00482_),
    .C(_00576_),
    .ZN(_00577_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06166_ (.I(_00519_),
    .Z(_00578_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06167_ (.I(\as2650.cycle[6] ),
    .Z(_00579_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06168_ (.I(_00579_),
    .Z(_00580_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06169_ (.I(_00580_),
    .Z(_00581_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06170_ (.I(_00581_),
    .Z(_00582_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06171_ (.I(_00582_),
    .Z(_00583_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06172_ (.I(_00583_),
    .Z(_00584_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06173_ (.A1(_00578_),
    .A2(_00584_),
    .ZN(_00585_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06174_ (.I(_00585_),
    .Z(_00586_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06175_ (.A1(_00548_),
    .A2(_00577_),
    .B(_00586_),
    .ZN(_00587_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06176_ (.I(_00468_),
    .Z(_00588_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06177_ (.I(_00588_),
    .Z(_00589_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06178_ (.I(_00476_),
    .Z(_00590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06179_ (.A1(_00590_),
    .A2(_05755_),
    .ZN(_00591_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06180_ (.A1(_00589_),
    .A2(_00591_),
    .ZN(_00592_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06181_ (.I(net6),
    .Z(_00593_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06182_ (.I(_00593_),
    .Z(_00594_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06183_ (.A1(_00594_),
    .A2(\as2650.cycle[1] ),
    .Z(_00595_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06184_ (.I(_00595_),
    .Z(_00596_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06185_ (.I(_00596_),
    .Z(_00597_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06186_ (.I(_00597_),
    .Z(_00598_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06187_ (.I(_00499_),
    .Z(_00599_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06188_ (.I(net3),
    .Z(_00600_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06189_ (.I(_00600_),
    .Z(_00601_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06190_ (.I(_00601_),
    .Z(_00602_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06191_ (.I(_00602_),
    .Z(_00603_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06192_ (.I(_00603_),
    .Z(_00604_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06193_ (.A1(_00599_),
    .A2(_00604_),
    .ZN(_00605_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06194_ (.A1(_00598_),
    .A2(_00605_),
    .ZN(_00606_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06195_ (.I(\as2650.cycle[9] ),
    .Z(_00607_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06196_ (.A1(_00593_),
    .A2(\as2650.cycle[1] ),
    .ZN(_00608_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06197_ (.I(_00608_),
    .Z(_00609_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06198_ (.I(_00609_),
    .Z(_00610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06199_ (.A1(_00593_),
    .A2(\as2650.cycle[10] ),
    .ZN(_00611_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06200_ (.I(net6),
    .Z(_00612_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06201_ (.I(_00612_),
    .Z(_00613_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06202_ (.A1(_00613_),
    .A2(\as2650.cycle[2] ),
    .ZN(_00614_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06203_ (.A1(_00611_),
    .A2(_00614_),
    .ZN(_00615_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06204_ (.I(_00615_),
    .Z(_00616_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06205_ (.A1(_00594_),
    .A2(\as2650.cycle[3] ),
    .Z(_00617_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06206_ (.I(_00617_),
    .Z(_00618_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06207_ (.A1(_05717_),
    .A2(_00616_),
    .A3(_00618_),
    .ZN(_00619_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06208_ (.A1(_00607_),
    .A2(_00610_),
    .A3(_00619_),
    .ZN(_00620_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06209_ (.A1(_00606_),
    .A2(_00620_),
    .ZN(_00621_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06210_ (.A1(_00486_),
    .A2(_05721_),
    .ZN(_00622_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06211_ (.A1(_00496_),
    .A2(_00622_),
    .ZN(_00623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06212_ (.I(_00623_),
    .Z(_00624_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06213_ (.I(_05754_),
    .Z(_00625_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06214_ (.I(_00625_),
    .Z(_00626_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06215_ (.I(_00626_),
    .Z(_00627_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _06216_ (.I(_00627_),
    .Z(_00628_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06217_ (.I(\as2650.addr_buff[7] ),
    .Z(_00629_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06218_ (.I(_00629_),
    .Z(_00630_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06219_ (.I(_00630_),
    .Z(_00631_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06220_ (.I(_00631_),
    .Z(_00632_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06221_ (.I(_00613_),
    .Z(_00633_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06222_ (.I(\as2650.cycle[10] ),
    .Z(_00634_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06223_ (.A1(_00633_),
    .A2(_00634_),
    .Z(_00635_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06224_ (.I(_00635_),
    .Z(_00636_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06225_ (.A1(_00595_),
    .A2(_00617_),
    .ZN(_00637_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06226_ (.I(_00637_),
    .Z(_00638_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06227_ (.A1(_00636_),
    .A2(_00638_),
    .ZN(_00639_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _06228_ (.A1(_00628_),
    .A2(_00506_),
    .A3(_00632_),
    .A4(_00639_),
    .ZN(_00640_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06229_ (.A1(_00621_),
    .A2(_00624_),
    .B1(_00640_),
    .B2(_00491_),
    .ZN(_00641_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06230_ (.I(\as2650.cycle[13] ),
    .Z(_00642_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06231_ (.A1(_00612_),
    .A2(_00642_),
    .ZN(_00643_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06232_ (.I(_00643_),
    .Z(_00644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06233_ (.A1(_00613_),
    .A2(\as2650.cycle[11] ),
    .ZN(_00645_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06234_ (.A1(_00644_),
    .A2(_00645_),
    .ZN(_00646_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06235_ (.I(_00646_),
    .Z(_00647_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06236_ (.A1(_00592_),
    .A2(_00641_),
    .A3(_00647_),
    .ZN(_00648_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06237_ (.A1(_00587_),
    .A2(_00648_),
    .ZN(_00649_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06238_ (.A1(_00575_),
    .A2(_00551_),
    .ZN(_00650_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06239_ (.A1(_00650_),
    .A2(_00647_),
    .ZN(_00651_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06240_ (.A1(_00610_),
    .A2(_00619_),
    .A3(_00651_),
    .ZN(_00652_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06241_ (.I(_00652_),
    .ZN(_00653_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06242_ (.I(_00645_),
    .Z(_00654_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06243_ (.I(_00484_),
    .Z(_00655_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _06244_ (.A1(net6),
    .A2(\as2650.cycle[13] ),
    .Z(_00656_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06245_ (.I(_00656_),
    .Z(_00657_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06246_ (.A1(_00655_),
    .A2(_00657_),
    .ZN(_00658_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06247_ (.A1(_00472_),
    .A2(_00658_),
    .ZN(_00659_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06248_ (.A1(_00612_),
    .A2(\as2650.cycle[5] ),
    .ZN(_00660_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06249_ (.I(_00660_),
    .Z(_00661_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06250_ (.I(\as2650.cycle[4] ),
    .Z(_00662_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06251_ (.A1(_00594_),
    .A2(_00662_),
    .ZN(_00663_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06252_ (.A1(_00545_),
    .A2(_00661_),
    .A3(_00663_),
    .ZN(_00664_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06253_ (.A1(_00659_),
    .A2(_00664_),
    .ZN(_00665_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06254_ (.A1(_00654_),
    .A2(_00665_),
    .ZN(_00666_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06255_ (.A1(net5),
    .A2(_00573_),
    .ZN(_00667_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06256_ (.I(_00667_),
    .Z(_00668_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06257_ (.I(_00522_),
    .Z(_00669_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06258_ (.I(_00568_),
    .Z(_00670_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06259_ (.A1(_00669_),
    .A2(_00670_),
    .ZN(_00671_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06260_ (.I(_00549_),
    .Z(_00672_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06261_ (.I(_00656_),
    .Z(_00673_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06262_ (.A1(_00672_),
    .A2(_00673_),
    .ZN(_00674_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06263_ (.I(_00674_),
    .Z(_00675_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06264_ (.A1(_00540_),
    .A2(_00675_),
    .ZN(_00676_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06265_ (.A1(_00671_),
    .A2(_00676_),
    .ZN(_00677_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06266_ (.I(_00509_),
    .Z(_00678_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06267_ (.I(_00521_),
    .Z(_00679_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06268_ (.I(_05748_),
    .Z(_00680_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06269_ (.A1(_00678_),
    .A2(_00679_),
    .A3(_00680_),
    .ZN(_00681_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06270_ (.I(_00681_),
    .Z(_00682_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06271_ (.I(_00527_),
    .Z(_00683_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _06272_ (.A1(_00678_),
    .A2(_00683_),
    .A3(_05844_),
    .Z(_00684_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06273_ (.I(_00684_),
    .Z(_00685_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06274_ (.A1(_00682_),
    .A2(_00685_),
    .ZN(_00686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06275_ (.I(_00524_),
    .Z(_00687_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06276_ (.I(\as2650.cycle[0] ),
    .Z(_00688_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06277_ (.I(net7),
    .ZN(_00689_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06278_ (.A1(_00689_),
    .A2(\as2650.last_intr ),
    .A3(net75),
    .ZN(_00690_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06279_ (.I(net72),
    .Z(_00691_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06280_ (.A1(_00688_),
    .A2(_00690_),
    .B(_00691_),
    .ZN(_00692_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06281_ (.A1(_05716_),
    .A2(_00692_),
    .ZN(_00693_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _06282_ (.A1(_00668_),
    .A2(_00677_),
    .B1(_00686_),
    .B2(_00687_),
    .C(_00693_),
    .ZN(_00694_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06283_ (.A1(_00633_),
    .A2(\as2650.cycle[7] ),
    .ZN(_00695_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06284_ (.I(\as2650.cycle[5] ),
    .Z(_00696_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06285_ (.A1(_00593_),
    .A2(_00696_),
    .Z(_00697_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06286_ (.I(_00697_),
    .Z(_00698_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06287_ (.I(_00698_),
    .Z(_00699_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06288_ (.I(_00657_),
    .Z(_00700_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06289_ (.A1(_00512_),
    .A2(_00700_),
    .ZN(_00701_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06290_ (.A1(_00594_),
    .A2(\as2650.cycle[12] ),
    .ZN(_00702_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06291_ (.A1(_00546_),
    .A2(_00701_),
    .A3(_00702_),
    .ZN(_00703_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06292_ (.A1(_05716_),
    .A2(_00699_),
    .A3(_00703_),
    .ZN(_00704_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06293_ (.I(_00528_),
    .Z(_00705_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _06294_ (.A1(_00705_),
    .A2(_00687_),
    .A3(_00681_),
    .A4(_00570_),
    .ZN(_00706_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06295_ (.A1(_00530_),
    .A2(_00706_),
    .ZN(_00707_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06296_ (.I(_00644_),
    .Z(_00708_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06297_ (.I(_00708_),
    .Z(_00709_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06298_ (.I(_00709_),
    .Z(_00710_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _06299_ (.A1(_00695_),
    .A2(_00704_),
    .B1(_00707_),
    .B2(_00710_),
    .ZN(_00711_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _06300_ (.A1(_00499_),
    .A2(_00666_),
    .B(_00694_),
    .C(_00711_),
    .ZN(_00712_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06301_ (.I(_00642_),
    .Z(_00713_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06302_ (.A1(_00653_),
    .A2(_00712_),
    .B(_00713_),
    .ZN(_00714_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06303_ (.A1(_00539_),
    .A2(_00649_),
    .A3(_00714_),
    .ZN(_00004_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06304_ (.I(_00510_),
    .Z(_00715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06305_ (.A1(_00526_),
    .A2(_00715_),
    .ZN(_00716_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06306_ (.I(_00716_),
    .Z(_00717_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06307_ (.I(_00717_),
    .Z(_00718_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06308_ (.I(_00718_),
    .Z(_00719_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06309_ (.A1(_00719_),
    .A2(_00491_),
    .ZN(_00720_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06310_ (.A1(\as2650.addr_buff[7] ),
    .A2(_00698_),
    .ZN(_00721_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06311_ (.A1(_05719_),
    .A2(_00467_),
    .A3(_00720_),
    .A4(_00721_),
    .ZN(_00722_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06312_ (.I(_00698_),
    .Z(_00723_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06313_ (.I(_00723_),
    .Z(_00724_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06314_ (.A1(_00679_),
    .A2(_00498_),
    .ZN(_00725_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06315_ (.I(_00725_),
    .Z(_00726_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06316_ (.A1(_00724_),
    .A2(_00726_),
    .ZN(_00727_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06317_ (.A1(_00504_),
    .A2(_00727_),
    .B(_00712_),
    .ZN(_00728_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06318_ (.A1(_00652_),
    .A2(_00728_),
    .ZN(_00729_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06319_ (.I(_00729_),
    .Z(_00730_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06320_ (.A1(_00701_),
    .A2(_00722_),
    .B1(_00730_),
    .B2(\as2650.cycle[12] ),
    .ZN(_00731_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06321_ (.I(_00731_),
    .ZN(_00003_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06322_ (.A1(_00540_),
    .A2(_00657_),
    .ZN(_00732_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06323_ (.I(_00732_),
    .Z(_00733_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06324_ (.I(_00733_),
    .Z(_00734_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06325_ (.I(_00599_),
    .Z(_00735_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06326_ (.I(_00735_),
    .Z(_00736_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06327_ (.A1(_00481_),
    .A2(_00472_),
    .ZN(_00737_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06328_ (.I(_00737_),
    .Z(_00738_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06329_ (.I(_00738_),
    .Z(_00739_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06330_ (.I(_00739_),
    .Z(_00740_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06331_ (.I(_00740_),
    .Z(_00741_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06332_ (.I(_00723_),
    .Z(_00742_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06333_ (.I(_00742_),
    .Z(_00743_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _06334_ (.A1(_00736_),
    .A2(_00741_),
    .A3(_00743_),
    .A4(_00663_),
    .ZN(_00744_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06335_ (.A1(_00547_),
    .A2(_00734_),
    .A3(_00744_),
    .ZN(_00745_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06336_ (.I(_00700_),
    .Z(_00746_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06337_ (.I(_00746_),
    .Z(_00747_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06338_ (.I(_00747_),
    .Z(_00748_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06339_ (.I(_00488_),
    .Z(_00749_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06340_ (.A1(_00499_),
    .A2(_00622_),
    .ZN(_00750_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06341_ (.A1(_00662_),
    .A2(_00749_),
    .A3(_00750_),
    .ZN(_00751_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06342_ (.A1(_00748_),
    .A2(_00751_),
    .ZN(_00752_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06343_ (.A1(\as2650.cycle[11] ),
    .A2(_00729_),
    .B1(_00752_),
    .B2(_00483_),
    .ZN(_00753_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06344_ (.A1(_00745_),
    .A2(_00753_),
    .ZN(_00002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06345_ (.A1(_00613_),
    .A2(\as2650.cycle[3] ),
    .ZN(_00754_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06346_ (.I(_00754_),
    .Z(_00755_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06347_ (.A1(_00597_),
    .A2(_00755_),
    .ZN(_00756_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06348_ (.A1(_00612_),
    .A2(\as2650.cycle[11] ),
    .Z(_00757_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06349_ (.I(_00757_),
    .Z(_00758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06350_ (.A1(_00623_),
    .A2(_00644_),
    .ZN(_00759_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06351_ (.I(_00759_),
    .Z(_00760_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06352_ (.A1(_00507_),
    .A2(_00758_),
    .A3(_00760_),
    .ZN(_00761_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06353_ (.A1(_00634_),
    .A2(_00730_),
    .B1(_00756_),
    .B2(_00761_),
    .ZN(_00762_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06354_ (.I(_00762_),
    .ZN(_00001_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06355_ (.I(\as2650.cycle[9] ),
    .ZN(_00763_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06356_ (.I(_00609_),
    .Z(_00764_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06357_ (.I(_00651_),
    .Z(_00765_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06358_ (.I(_00618_),
    .Z(_00766_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06359_ (.I(_00633_),
    .Z(_00767_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06360_ (.I(\as2650.cycle[2] ),
    .Z(_00768_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06361_ (.I(_00611_),
    .Z(_00769_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06362_ (.A1(_00767_),
    .A2(_00768_),
    .A3(_00769_),
    .ZN(_00770_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06363_ (.A1(_00736_),
    .A2(_00766_),
    .A3(_00770_),
    .ZN(_00771_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06364_ (.A1(_00764_),
    .A2(_00765_),
    .A3(_00771_),
    .ZN(_00772_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06365_ (.A1(_00763_),
    .A2(_00728_),
    .B(_00772_),
    .ZN(_00013_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06366_ (.I(_00736_),
    .Z(_00773_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06367_ (.A1(_00691_),
    .A2(_00690_),
    .ZN(_00774_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06368_ (.I(_00749_),
    .Z(_00775_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06369_ (.I(_00775_),
    .Z(_00776_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06370_ (.I(_00776_),
    .Z(_00777_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06371_ (.A1(_00767_),
    .A2(_00777_),
    .ZN(_00778_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06372_ (.I(\as2650.cycle[8] ),
    .Z(_00779_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06373_ (.I(_00779_),
    .Z(_00780_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06374_ (.I(_00780_),
    .Z(_00781_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06375_ (.I(_00781_),
    .Z(_00782_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06376_ (.I(_00782_),
    .Z(_00783_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06377_ (.I(_00783_),
    .Z(_00784_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06378_ (.A1(_00688_),
    .A2(_00774_),
    .B1(_00778_),
    .B2(_00784_),
    .ZN(_00785_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06379_ (.A1(_00773_),
    .A2(_00785_),
    .ZN(_00012_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06380_ (.I(_00660_),
    .Z(_00786_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06381_ (.I(_00786_),
    .Z(_00787_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06382_ (.A1(_00787_),
    .A2(_00701_),
    .ZN(_00788_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06383_ (.A1(_00736_),
    .A2(_00702_),
    .A3(_00788_),
    .ZN(_00789_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06384_ (.A1(\as2650.cycle[7] ),
    .A2(_00730_),
    .B1(_00789_),
    .B2(_00547_),
    .ZN(_00790_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06385_ (.I(_00790_),
    .ZN(_00011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06386_ (.I(_00580_),
    .Z(_00791_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06387_ (.I(_00791_),
    .Z(_00792_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06388_ (.I(_00792_),
    .Z(_00793_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06389_ (.I(_00793_),
    .Z(_00794_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06390_ (.I(_00794_),
    .Z(_00795_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06391_ (.I(_00795_),
    .Z(_00796_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06392_ (.I(_00779_),
    .ZN(_00797_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06393_ (.I(_00797_),
    .Z(_00798_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06394_ (.I(_00798_),
    .Z(_00799_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06395_ (.I(_00520_),
    .Z(_00800_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06396_ (.A1(_00799_),
    .A2(_00800_),
    .ZN(_00801_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06397_ (.I(_00801_),
    .Z(_00802_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06398_ (.A1(_00796_),
    .A2(_00693_),
    .B1(_00802_),
    .B2(_00767_),
    .ZN(_00803_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06399_ (.I(_00803_),
    .ZN(_00010_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _06400_ (.I(_00696_),
    .ZN(_00804_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06401_ (.I(_00804_),
    .Z(_00805_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06402_ (.I(_00805_),
    .Z(_00806_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06403_ (.I(_00622_),
    .Z(_00807_));
 gf180mcu_fd_sc_mcu7t5v0__or2_4 _06404_ (.A1(\as2650.ins_reg[2] ),
    .A2(\as2650.ins_reg[3] ),
    .Z(_00808_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06405_ (.I(_00808_),
    .Z(_00809_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06406_ (.I(_00809_),
    .Z(_00810_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06407_ (.I(_00810_),
    .Z(_00811_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06408_ (.I(_00811_),
    .Z(_00812_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06409_ (.I(_00812_),
    .Z(_00813_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06410_ (.A1(_05754_),
    .A2(_00477_),
    .A3(_00813_),
    .ZN(_00814_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06411_ (.I(_00814_),
    .Z(_00815_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06412_ (.A1(_05842_),
    .A2(_05747_),
    .ZN(_00816_));
 gf180mcu_fd_sc_mcu7t5v0__and2_4 _06413_ (.A1(_00680_),
    .A2(_00816_),
    .Z(_00817_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06414_ (.A1(_00585_),
    .A2(_00807_),
    .A3(_00815_),
    .A4(_00817_),
    .ZN(_00818_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06415_ (.I(_00557_),
    .Z(_00819_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06416_ (.I(_00819_),
    .Z(_00820_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06417_ (.A1(_00494_),
    .A2(_00820_),
    .ZN(_00821_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _06418_ (.A1(_00521_),
    .A2(_00591_),
    .A3(_00821_),
    .Z(_00822_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06419_ (.A1(_00525_),
    .A2(_00822_),
    .ZN(_00823_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06420_ (.A1(_00813_),
    .A2(_00823_),
    .ZN(_00824_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06421_ (.I(_00626_),
    .Z(_00825_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06422_ (.I(_00825_),
    .Z(_00826_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06423_ (.I(_00826_),
    .Z(_00827_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06424_ (.I(_00678_),
    .Z(_00828_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06425_ (.I(_00828_),
    .Z(_00829_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06426_ (.I(_00829_),
    .Z(_00830_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06427_ (.I(_00830_),
    .Z(_00831_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06428_ (.I(_00464_),
    .Z(_00832_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06429_ (.I(_00832_),
    .Z(_00833_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06430_ (.I(_00833_),
    .Z(_00834_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06431_ (.A1(_00831_),
    .A2(_00834_),
    .ZN(_00835_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06432_ (.I(_00549_),
    .Z(_00836_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06433_ (.I(_00836_),
    .Z(_00837_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06434_ (.I(_00837_),
    .Z(_00838_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06435_ (.I(_00838_),
    .Z(_00839_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06436_ (.I(_00839_),
    .Z(_00840_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06437_ (.A1(_00827_),
    .A2(_00835_),
    .B(_00735_),
    .C(_00840_),
    .ZN(_00841_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _06438_ (.A1(_00818_),
    .A2(_00824_),
    .B1(_00841_),
    .B2(_00748_),
    .ZN(_00842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06439_ (.A1(_00713_),
    .A2(_00505_),
    .ZN(_00843_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _06440_ (.A1(_00806_),
    .A2(_00728_),
    .B1(_00842_),
    .B2(_00496_),
    .C(_00843_),
    .ZN(_00009_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _06441_ (.I(_00662_),
    .ZN(_00844_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06442_ (.I(_00578_),
    .Z(_00845_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06443_ (.I(_00845_),
    .Z(_00846_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06444_ (.I(net3),
    .Z(_00847_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06445_ (.I(_00847_),
    .Z(_00848_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06446_ (.I(_00848_),
    .Z(_00849_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06447_ (.I(_00849_),
    .Z(_00850_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06448_ (.I(_00850_),
    .Z(_00851_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06449_ (.I(_00851_),
    .Z(_00852_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06450_ (.I(_00717_),
    .Z(_00853_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06451_ (.I(_00853_),
    .Z(_00854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06452_ (.I(_00489_),
    .Z(_00855_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06453_ (.I(_00855_),
    .Z(_00856_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06454_ (.I(_00710_),
    .Z(_00857_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06455_ (.I(_00700_),
    .Z(_00858_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06456_ (.A1(_00526_),
    .A2(_00858_),
    .ZN(_00859_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06457_ (.I(_00859_),
    .Z(_00860_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06458_ (.I(_00466_),
    .Z(_00861_));
 gf180mcu_fd_sc_mcu7t5v0__oai33_4 _06459_ (.A1(_00854_),
    .A2(_00856_),
    .A3(_00857_),
    .B1(_00860_),
    .B2(_00720_),
    .B3(_00861_),
    .ZN(_00862_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06460_ (.A1(_00846_),
    .A2(_00852_),
    .A3(_00862_),
    .ZN(_00863_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06461_ (.A1(_00737_),
    .A2(_00656_),
    .ZN(_00864_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06462_ (.I(_00596_),
    .Z(_00865_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06463_ (.I(_00865_),
    .Z(_00866_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _06464_ (.A1(_05718_),
    .A2(_00632_),
    .A3(_00639_),
    .B1(_00620_),
    .B2(_00628_),
    .ZN(_00867_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06465_ (.A1(_00866_),
    .A2(_00605_),
    .B(_00867_),
    .ZN(_00868_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06466_ (.A1(_00477_),
    .A2(_00868_),
    .ZN(_00869_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06467_ (.A1(_00722_),
    .A2(_00864_),
    .B1(_00869_),
    .B2(_00765_),
    .ZN(_00870_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06468_ (.A1(_00844_),
    .A2(_00728_),
    .B(_00863_),
    .C(_00870_),
    .ZN(_00008_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06469_ (.A1(_00586_),
    .A2(_00807_),
    .A3(_00835_),
    .ZN(_00871_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06470_ (.A1(\as2650.cycle[3] ),
    .A2(_00730_),
    .B1(_00871_),
    .B2(_00576_),
    .ZN(_00872_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06471_ (.I(_00872_),
    .ZN(_00007_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06472_ (.A1(_05754_),
    .A2(_00489_),
    .ZN(_00873_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06473_ (.I(_00470_),
    .Z(_00874_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06474_ (.I(_00874_),
    .Z(_00875_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06475_ (.I(_00875_),
    .Z(_00876_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06476_ (.I(_00876_),
    .Z(_00877_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06477_ (.A1(_00831_),
    .A2(_00877_),
    .A3(_00586_),
    .ZN(_00878_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06478_ (.A1(\as2650.cycle[1] ),
    .A2(_00729_),
    .B1(_00873_),
    .B2(_00878_),
    .ZN(_00879_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06479_ (.I(_00879_),
    .ZN(_00005_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06480_ (.A1(_00768_),
    .A2(_00729_),
    .ZN(_00880_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06481_ (.A1(_00852_),
    .A2(_00866_),
    .A3(_00761_),
    .ZN(_00881_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06482_ (.I(_00578_),
    .Z(_00882_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06483_ (.I(_00882_),
    .Z(_00883_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06484_ (.A1(_00608_),
    .A2(_00754_),
    .ZN(_00884_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06485_ (.A1(_00769_),
    .A2(_00884_),
    .ZN(_00885_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _06486_ (.A1(_00883_),
    .A2(_00632_),
    .A3(_00885_),
    .A4(_00765_),
    .ZN(_00886_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06487_ (.A1(_00880_),
    .A2(_00881_),
    .A3(_00886_),
    .ZN(_00006_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06488_ (.A1(_05751_),
    .A2(_00459_),
    .Z(_00887_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06489_ (.I(_00887_),
    .Z(_00888_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _06490_ (.A1(\as2650.addr_buff[7] ),
    .A2(_00660_),
    .Z(_00889_));
 gf180mcu_fd_sc_mcu7t5v0__oai33_1 _06491_ (.A1(_00888_),
    .A2(_00741_),
    .A3(_00586_),
    .B1(_00748_),
    .B2(_00889_),
    .B3(_00735_),
    .ZN(_00890_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06492_ (.A1(_00854_),
    .A2(_00547_),
    .A3(_00890_),
    .ZN(_00891_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06493_ (.I(_00503_),
    .Z(_00892_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06494_ (.I(_00570_),
    .Z(_00893_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06495_ (.I(_00655_),
    .Z(_00894_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06496_ (.I(_00709_),
    .Z(_00895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06497_ (.A1(_00468_),
    .A2(_00501_),
    .ZN(_00896_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06498_ (.I(_00896_),
    .Z(_00897_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06499_ (.A1(_00897_),
    .A2(_00682_),
    .ZN(_00898_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06500_ (.A1(_00894_),
    .A2(_00895_),
    .A3(_00898_),
    .ZN(_00899_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _06501_ (.A1(_00892_),
    .A2(_00687_),
    .A3(_00893_),
    .A4(_00899_),
    .Z(_00900_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06502_ (.I(_00494_),
    .Z(_00901_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06503_ (.I(_00901_),
    .Z(_00902_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06504_ (.I(_00560_),
    .Z(_00903_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06505_ (.A1(_00902_),
    .A2(_00478_),
    .A3(_00903_),
    .ZN(_00904_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06506_ (.I(_05721_),
    .Z(_00905_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06507_ (.I(_00905_),
    .Z(_00906_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06508_ (.A1(_00906_),
    .A2(_00534_),
    .ZN(_00907_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06509_ (.A1(_00856_),
    .A2(_00904_),
    .A3(_00907_),
    .ZN(_00908_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06510_ (.I(_05717_),
    .Z(_00909_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06511_ (.A1(_00688_),
    .A2(_00693_),
    .B(_00908_),
    .C(_00909_),
    .ZN(_00910_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _06512_ (.A1(_00826_),
    .A2(_00805_),
    .A3(_00856_),
    .B1(_00751_),
    .B2(_00483_),
    .ZN(_00911_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06513_ (.I(_00486_),
    .Z(_00912_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06514_ (.I(_00912_),
    .Z(_00913_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06515_ (.I(_00913_),
    .Z(_00914_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06516_ (.A1(\as2650.cycle[5] ),
    .A2(\as2650.cycle[4] ),
    .ZN(_00915_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06517_ (.I(_00915_),
    .Z(_00916_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06518_ (.I(_00916_),
    .Z(_00917_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06519_ (.I(_00581_),
    .Z(_00918_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06520_ (.I(_00918_),
    .Z(_00919_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _06521_ (.A1(_00688_),
    .A2(_00713_),
    .A3(_00919_),
    .A4(\as2650.cycle[11] ),
    .ZN(_00920_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06522_ (.A1(_00607_),
    .A2(\as2650.cycle[12] ),
    .A3(\as2650.cycle[7] ),
    .ZN(_00921_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _06523_ (.A1(\as2650.cycle[1] ),
    .A2(\as2650.cycle[3] ),
    .A3(_00634_),
    .A4(_00768_),
    .ZN(_00922_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _06524_ (.A1(_00917_),
    .A2(_00920_),
    .A3(_00921_),
    .A4(_00922_),
    .Z(_00923_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _06525_ (.A1(_00914_),
    .A2(_00495_),
    .B(_00800_),
    .C(_00923_),
    .ZN(_00924_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06526_ (.A1(_00658_),
    .A2(_00911_),
    .B(_00924_),
    .ZN(_00925_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06527_ (.A1(_00530_),
    .A2(_00857_),
    .B(_00910_),
    .C(_00925_),
    .ZN(_00926_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06528_ (.I(_00787_),
    .Z(_00927_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06529_ (.I(_00927_),
    .Z(_00928_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _06530_ (.A1(_00735_),
    .A2(_00892_),
    .A3(_00928_),
    .A4(_00726_),
    .ZN(_00929_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _06531_ (.A1(_05719_),
    .A2(_00743_),
    .A3(_00695_),
    .A4(_00703_),
    .ZN(_00930_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _06532_ (.A1(_00900_),
    .A2(_00926_),
    .A3(_00929_),
    .A4(_00930_),
    .ZN(_00931_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06533_ (.A1(_00659_),
    .A2(_00664_),
    .B(_00760_),
    .ZN(_00932_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _06534_ (.A1(_00605_),
    .A2(_00862_),
    .B1(_00932_),
    .B2(_00758_),
    .ZN(_00933_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06535_ (.A1(_00490_),
    .A2(_00561_),
    .ZN(_00934_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06536_ (.A1(_00476_),
    .A2(_05753_),
    .A3(_05748_),
    .ZN(_00935_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06537_ (.I(_05782_),
    .Z(_00936_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06538_ (.A1(_00936_),
    .A2(_00560_),
    .ZN(_00937_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06539_ (.A1(_00935_),
    .A2(_00937_),
    .ZN(_00938_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06540_ (.I(_00938_),
    .Z(_00939_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06541_ (.A1(_00821_),
    .A2(_00935_),
    .ZN(_00940_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06542_ (.I(_00940_),
    .Z(_00941_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06543_ (.I(_00941_),
    .Z(_00942_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06544_ (.I(_05744_),
    .Z(_00943_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06545_ (.A1(_00943_),
    .A2(_00566_),
    .A3(_00937_),
    .ZN(_00944_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06546_ (.A1(_00939_),
    .A2(_00942_),
    .A3(_00944_),
    .ZN(_00945_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06547_ (.I(_05773_),
    .Z(_00946_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06548_ (.I(_00946_),
    .Z(_00947_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06549_ (.I(_00555_),
    .Z(_00948_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06550_ (.I(_00903_),
    .Z(_00949_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _06551_ (.A1(_00947_),
    .A2(_00948_),
    .A3(_00949_),
    .A4(_00572_),
    .ZN(_00950_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06552_ (.A1(_00624_),
    .A2(_00823_),
    .ZN(_00951_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06553_ (.A1(_00934_),
    .A2(_00945_),
    .B(_00950_),
    .C(_00951_),
    .ZN(_00952_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06554_ (.I(_00522_),
    .Z(_00953_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06555_ (.A1(_00575_),
    .A2(_00953_),
    .ZN(_00954_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06556_ (.A1(_00680_),
    .A2(_00816_),
    .ZN(_00955_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06557_ (.I(_00955_),
    .Z(_00956_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _06558_ (.A1(_00831_),
    .A2(_05719_),
    .A3(_00954_),
    .A4(_00956_),
    .ZN(_00957_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _06559_ (.A1(_00750_),
    .A2(_00815_),
    .A3(_00956_),
    .A4(_00904_),
    .ZN(_00958_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06560_ (.I(_00953_),
    .Z(_00959_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06561_ (.I(_00959_),
    .Z(_00960_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06562_ (.I(_00567_),
    .Z(_00961_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _06563_ (.A1(_00678_),
    .A2(_00566_),
    .A3(_00961_),
    .Z(_00962_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06564_ (.I(_00962_),
    .Z(_00963_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06565_ (.A1(_00527_),
    .A2(_05749_),
    .ZN(_00964_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06566_ (.A1(_00946_),
    .A2(_00903_),
    .A3(_00964_),
    .ZN(_00965_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06567_ (.I(_00574_),
    .Z(_00966_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06568_ (.I(_00966_),
    .Z(_00967_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06569_ (.I(_00967_),
    .Z(_00968_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06570_ (.I(_00968_),
    .Z(_00969_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _06571_ (.A1(_00800_),
    .A2(_00963_),
    .B1(_00965_),
    .B2(_00969_),
    .ZN(_00970_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06572_ (.I(_05736_),
    .Z(_00971_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06573_ (.I(_05728_),
    .Z(_00972_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06574_ (.A1(_00972_),
    .A2(_00812_),
    .A3(_00935_),
    .ZN(_00973_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06575_ (.I(_00973_),
    .Z(_00974_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06576_ (.A1(_00971_),
    .A2(_00974_),
    .ZN(_00975_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06577_ (.A1(_00565_),
    .A2(_00975_),
    .ZN(_00976_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06578_ (.A1(_00960_),
    .A2(_00970_),
    .B(_00976_),
    .ZN(_00977_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06579_ (.I(_00561_),
    .Z(_00978_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06580_ (.A1(_00837_),
    .A2(_00978_),
    .ZN(_00979_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06581_ (.I(_00820_),
    .Z(_00980_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06582_ (.A1(_05763_),
    .A2(_00948_),
    .A3(_00980_),
    .ZN(_00981_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06583_ (.I(_00981_),
    .Z(_00982_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06584_ (.I(_00982_),
    .Z(_00983_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06585_ (.I(_00983_),
    .Z(_00984_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06586_ (.A1(_00856_),
    .A2(_00984_),
    .ZN(_00985_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06587_ (.A1(_00687_),
    .A2(_00686_),
    .B1(_00979_),
    .B2(_00668_),
    .C(_00985_),
    .ZN(_00986_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06588_ (.A1(_00496_),
    .A2(_00958_),
    .B(_00977_),
    .C(_00986_),
    .ZN(_00987_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _06589_ (.A1(_00952_),
    .A2(_00957_),
    .A3(_00987_),
    .B(_00538_),
    .ZN(_00988_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _06590_ (.A1(_00891_),
    .A2(_00931_),
    .A3(_00933_),
    .A4(_00988_),
    .ZN(_00000_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06591_ (.I(net28),
    .ZN(net15));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06592_ (.I(_00936_),
    .Z(_00989_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06593_ (.A1(_05781_),
    .A2(_00475_),
    .ZN(_00990_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _06594_ (.I(\as2650.cycle[6] ),
    .ZN(_00991_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06595_ (.A1(\as2650.cycle[8] ),
    .A2(_00991_),
    .ZN(_00992_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06596_ (.A1(_00667_),
    .A2(_00992_),
    .ZN(_00993_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06597_ (.A1(_00990_),
    .A2(_00993_),
    .ZN(_00994_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06598_ (.A1(_00962_),
    .A2(_00684_),
    .ZN(_00995_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06599_ (.A1(_00959_),
    .A2(_00995_),
    .ZN(_00996_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06600_ (.I(_05756_),
    .Z(_00997_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06601_ (.A1(_00997_),
    .A2(_00544_),
    .ZN(_00998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06602_ (.A1(_00996_),
    .A2(_00998_),
    .ZN(_00999_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06603_ (.A1(_05780_),
    .A2(_00901_),
    .ZN(_01000_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06604_ (.A1(\as2650.cycle[8] ),
    .A2(_00520_),
    .ZN(_01001_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06605_ (.I(_01001_),
    .Z(_01002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06606_ (.A1(_00991_),
    .A2(_00522_),
    .ZN(_01003_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06607_ (.A1(_00896_),
    .A2(_01003_),
    .ZN(_01004_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _06608_ (.A1(_00673_),
    .A2(_01000_),
    .A3(_01002_),
    .A4(_01004_),
    .Z(_01005_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06609_ (.I(_01005_),
    .Z(_01006_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06610_ (.I(_05780_),
    .Z(_01007_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06611_ (.I(_01007_),
    .Z(_01008_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06612_ (.I(\as2650.idx_ctrl[1] ),
    .Z(_01009_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06613_ (.A1(_01009_),
    .A2(\as2650.idx_ctrl[0] ),
    .ZN(_01010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06614_ (.A1(_00474_),
    .A2(_01010_),
    .ZN(_01011_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06615_ (.I(_01011_),
    .Z(_01012_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06616_ (.A1(_00590_),
    .A2(_00588_),
    .A3(_05742_),
    .ZN(_01013_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _06617_ (.A1(_00804_),
    .A2(_00980_),
    .A3(_01012_),
    .A4(_01013_),
    .Z(_01014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _06618_ (.A1(_00551_),
    .A2(_01002_),
    .ZN(_01015_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06619_ (.I(_00991_),
    .Z(_01016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06620_ (.A1(_01016_),
    .A2(_00644_),
    .ZN(_01017_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06621_ (.I(_01017_),
    .Z(_01018_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06622_ (.A1(_01008_),
    .A2(_01014_),
    .A3(_01015_),
    .A4(_01018_),
    .ZN(_01019_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _06623_ (.A1(_00994_),
    .A2(_00999_),
    .B(_01006_),
    .C(_01019_),
    .ZN(_01020_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06624_ (.I(_01000_),
    .Z(_01021_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06625_ (.A1(_00672_),
    .A2(_00993_),
    .ZN(_01022_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06626_ (.A1(_00814_),
    .A2(_01021_),
    .A3(_01022_),
    .ZN(_01023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06627_ (.I(_01023_),
    .Z(_01024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06628_ (.I(_01010_),
    .Z(_01025_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06629_ (.I(_01025_),
    .Z(_01026_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06630_ (.A1(_00550_),
    .A2(_00916_),
    .A3(_01002_),
    .ZN(_01027_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06631_ (.A1(_00615_),
    .A2(_01026_),
    .A3(_01017_),
    .A4(_01027_),
    .ZN(_01028_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06632_ (.A1(_00763_),
    .A2(_00884_),
    .A3(_00757_),
    .ZN(_01029_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06633_ (.A1(_01021_),
    .A2(_01028_),
    .A3(_01029_),
    .ZN(_01030_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06634_ (.A1(_00580_),
    .A2(_00646_),
    .ZN(_01031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06635_ (.A1(_00885_),
    .A2(_01031_),
    .ZN(_01032_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06636_ (.I(_00696_),
    .Z(_01033_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _06637_ (.A1(_01033_),
    .A2(_00662_),
    .A3(_01015_),
    .ZN(_01034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06638_ (.I(\as2650.addr_buff[6] ),
    .Z(_01035_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06639_ (.I(\as2650.addr_buff[5] ),
    .Z(_01036_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06640_ (.A1(_01035_),
    .A2(_01036_),
    .ZN(_01037_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06641_ (.A1(\as2650.addr_buff[7] ),
    .A2(_01037_),
    .ZN(_01038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06642_ (.A1(_01034_),
    .A2(_01038_),
    .ZN(_01039_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06643_ (.A1(_00990_),
    .A2(_01032_),
    .A3(_01039_),
    .ZN(_01040_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06644_ (.I(_01040_),
    .ZN(_01041_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06645_ (.A1(_01024_),
    .A2(_01030_),
    .A3(_01041_),
    .Z(_01042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06646_ (.A1(_01020_),
    .A2(_01042_),
    .ZN(_01043_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06647_ (.I(_01043_),
    .Z(_01044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06648_ (.A1(_00989_),
    .A2(_01044_),
    .ZN(_01045_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06649_ (.I(_01045_),
    .Z(_01046_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06650_ (.I(_01019_),
    .Z(_01047_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06651_ (.I(\as2650.idx_ctrl[1] ),
    .ZN(_01048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06652_ (.I(\as2650.idx_ctrl[0] ),
    .Z(_01049_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _06653_ (.A1(_01048_),
    .A2(_01049_),
    .A3(_05841_),
    .Z(_01050_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06654_ (.I(_01050_),
    .Z(_01051_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06655_ (.I(_05830_),
    .Z(_01052_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06656_ (.I(_01052_),
    .Z(_01053_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06657_ (.I(_01053_),
    .Z(_01054_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06658_ (.I(_01024_),
    .Z(_01055_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _06659_ (.A1(_00885_),
    .A2(_01031_),
    .Z(_01056_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _06660_ (.A1(_01021_),
    .A2(_01034_),
    .A3(_01038_),
    .A4(_01056_),
    .ZN(_01057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06661_ (.I(_01057_),
    .Z(_01058_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06662_ (.I(_01023_),
    .Z(_01059_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06663_ (.I(_00993_),
    .Z(_01060_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06664_ (.I(_00569_),
    .Z(_01061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06665_ (.A1(_00669_),
    .A2(_01061_),
    .ZN(_01062_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06666_ (.I(_01062_),
    .Z(_01063_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06667_ (.A1(_00990_),
    .A2(_01060_),
    .A3(_01063_),
    .ZN(_01064_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06668_ (.I(net50),
    .Z(_01065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06669_ (.I(_05785_),
    .Z(_01066_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06670_ (.I(_01066_),
    .Z(_01067_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06671_ (.A1(net50),
    .A2(net78),
    .ZN(_01068_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06672_ (.I(_01068_),
    .Z(_01069_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06673_ (.A1(_01065_),
    .A2(_01067_),
    .B(_01069_),
    .ZN(_01070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06674_ (.A1(_01064_),
    .A2(_01070_),
    .ZN(_01071_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06675_ (.I(_00442_),
    .Z(_01072_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06676_ (.I(_01072_),
    .ZN(_01073_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06677_ (.A1(_00669_),
    .A2(_00568_),
    .A3(_00994_),
    .ZN(_01074_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06678_ (.I(_01074_),
    .Z(_01075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06679_ (.I(_01075_),
    .Z(_01076_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06680_ (.I(_01074_),
    .Z(_01077_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06681_ (.I(net8),
    .Z(_01078_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06682_ (.I(_01078_),
    .Z(_01079_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06683_ (.I(_01079_),
    .Z(_01080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06684_ (.A1(_01080_),
    .A2(_01005_),
    .ZN(_01081_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06685_ (.A1(_00455_),
    .A2(_01006_),
    .B(_01077_),
    .C(_01081_),
    .ZN(_01082_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06686_ (.A1(_00669_),
    .A2(_00569_),
    .A3(_00994_),
    .ZN(_01083_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06687_ (.I(_01083_),
    .Z(_01084_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06688_ (.A1(_01073_),
    .A2(_01076_),
    .B(_01082_),
    .C(_01084_),
    .ZN(_01085_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06689_ (.A1(_01059_),
    .A2(_01071_),
    .A3(_01085_),
    .ZN(_01086_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06690_ (.A1(_01054_),
    .A2(_01055_),
    .B(_01058_),
    .C(_01086_),
    .ZN(_01087_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _06691_ (.A1(_00629_),
    .A2(_01037_),
    .Z(_01088_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _06692_ (.A1(_00990_),
    .A2(_01027_),
    .A3(_01088_),
    .A4(_01032_),
    .ZN(_01089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06693_ (.I(_01089_),
    .Z(_01090_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _06694_ (.I(\as2650.addr_buff[6] ),
    .ZN(_01091_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06695_ (.A1(_01091_),
    .A2(\as2650.addr_buff[5] ),
    .Z(_01092_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06696_ (.A1(_05841_),
    .A2(_01092_),
    .Z(_01093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06697_ (.I(_01093_),
    .Z(_01094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06698_ (.A1(_01090_),
    .A2(_01094_),
    .ZN(_01095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06699_ (.A1(_01087_),
    .A2(_01095_),
    .ZN(_01096_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06700_ (.I(_01030_),
    .Z(_01097_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06701_ (.I0(_01051_),
    .I1(_01096_),
    .S(_01097_),
    .Z(_01098_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06702_ (.I(\as2650.holding_reg[0] ),
    .Z(_01099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06703_ (.A1(_00445_),
    .A2(_00557_),
    .ZN(_01100_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _06704_ (.A1(_05773_),
    .A2(_05832_),
    .B1(_05831_),
    .B2(_05859_),
    .ZN(_01101_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06705_ (.A1(_01009_),
    .A2(_01049_),
    .Z(_01102_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06706_ (.I(_01102_),
    .Z(_01103_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06707_ (.A1(_05762_),
    .A2(_01103_),
    .B(_01052_),
    .ZN(_01104_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06708_ (.I(_00808_),
    .Z(_01105_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _06709_ (.A1(_01101_),
    .A2(_01103_),
    .B(_01104_),
    .C(_01105_),
    .ZN(_01106_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06710_ (.A1(_01099_),
    .A2(_01100_),
    .A3(_01106_),
    .ZN(_01107_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06711_ (.I(_00590_),
    .Z(_01108_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _06712_ (.A1(_01108_),
    .A2(_00589_),
    .A3(_00997_),
    .ZN(_01109_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06713_ (.I(_00683_),
    .Z(_01110_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06714_ (.A1(_01110_),
    .A2(_00588_),
    .A3(_05756_),
    .ZN(_01111_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06715_ (.I(_01111_),
    .Z(_01112_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06716_ (.A1(\as2650.holding_reg[0] ),
    .A2(_01105_),
    .Z(_01113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06717_ (.A1(\as2650.holding_reg[0] ),
    .A2(_00809_),
    .ZN(_01114_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06718_ (.A1(_00444_),
    .A2(_01105_),
    .B(_01114_),
    .ZN(_01115_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06719_ (.A1(_01106_),
    .A2(_01113_),
    .B(_01115_),
    .ZN(_01116_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06720_ (.I(_05744_),
    .Z(_01117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06721_ (.I(_05742_),
    .Z(_01118_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06722_ (.A1(_00683_),
    .A2(_00588_),
    .A3(_01118_),
    .ZN(_01119_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06723_ (.A1(_01117_),
    .A2(_00961_),
    .A3(_01119_),
    .ZN(_01120_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06724_ (.I(_01120_),
    .Z(_01121_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _06725_ (.A1(_01107_),
    .A2(_01109_),
    .B1(_01112_),
    .B2(_01116_),
    .C(_01121_),
    .ZN(_01122_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06726_ (.A1(_01099_),
    .A2(_01100_),
    .A3(_01106_),
    .Z(_01123_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06727_ (.A1(_01123_),
    .A2(_01116_),
    .Z(_01124_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06728_ (.I(_01124_),
    .Z(_01125_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06729_ (.A1(_01110_),
    .A2(_00943_),
    .ZN(_01126_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06730_ (.I(_01126_),
    .Z(_01127_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06731_ (.A1(_01069_),
    .A2(_01125_),
    .B(_01127_),
    .ZN(_01128_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06732_ (.A1(_01069_),
    .A2(_01125_),
    .B(_01128_),
    .ZN(_01129_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06733_ (.I(_01119_),
    .Z(_01130_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06734_ (.I(_01130_),
    .Z(_01131_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06735_ (.I(net78),
    .ZN(_01132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06736_ (.A1(net50),
    .A2(_01132_),
    .ZN(_01133_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06737_ (.A1(_01124_),
    .A2(_01133_),
    .Z(_01134_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06738_ (.A1(_00590_),
    .A2(_00589_),
    .A3(_00997_),
    .ZN(_01135_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06739_ (.A1(_01124_),
    .A2(_01133_),
    .B(_01135_),
    .ZN(_01136_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _06740_ (.A1(_01131_),
    .A2(_01125_),
    .B1(_01134_),
    .B2(_01136_),
    .ZN(_01137_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06741_ (.I(_01120_),
    .Z(_01138_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _06742_ (.A1(_01122_),
    .A2(_01129_),
    .A3(_01137_),
    .B1(_01115_),
    .B2(_01138_),
    .ZN(_01139_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06743_ (.A1(_01047_),
    .A2(net82),
    .ZN(_01140_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06744_ (.A1(_01047_),
    .A2(_01098_),
    .B(_01140_),
    .ZN(_01141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06745_ (.I(_01054_),
    .Z(_01142_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06746_ (.I0(\as2650.r123[0][0] ),
    .I1(\as2650.r123_2[0][0] ),
    .S(_05774_),
    .Z(_01143_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06747_ (.I(_01143_),
    .Z(_01144_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06748_ (.I(_01144_),
    .Z(_01145_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06749_ (.I(_01145_),
    .Z(_01146_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06750_ (.I(_05781_),
    .Z(_01147_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06751_ (.I(_01022_),
    .Z(_01148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06752_ (.A1(_01147_),
    .A2(_01148_),
    .ZN(_01149_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06753_ (.A1(_00978_),
    .A2(_01149_),
    .ZN(_01150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06754_ (.I(_01150_),
    .Z(_01151_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06755_ (.A1(_01142_),
    .A2(_01146_),
    .A3(_01151_),
    .ZN(_01152_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _06756_ (.A1(_00989_),
    .A2(_01044_),
    .B(_01151_),
    .C(_00506_),
    .ZN(_01153_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06757_ (.I(_01153_),
    .Z(_01154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06758_ (.A1(\as2650.r123[1][0] ),
    .A2(_01154_),
    .ZN(_01155_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06759_ (.A1(_01046_),
    .A2(_01141_),
    .B(_01152_),
    .C(_01155_),
    .ZN(_00014_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06760_ (.I(_01045_),
    .Z(_01156_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06761_ (.I(_01135_),
    .Z(_01157_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06762_ (.A1(_01123_),
    .A2(_01116_),
    .B(_01133_),
    .ZN(_01158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06763_ (.A1(\as2650.holding_reg[1] ),
    .A2(_00808_),
    .ZN(_01159_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06764_ (.A1(_00431_),
    .A2(_00809_),
    .B(_01159_),
    .ZN(_01160_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06765_ (.I(\as2650.holding_reg[1] ),
    .ZN(_01161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06766_ (.A1(_05772_),
    .A2(_05826_),
    .B1(_05825_),
    .B2(_05859_),
    .ZN(_01162_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06767_ (.A1(_01162_),
    .A2(_01102_),
    .Z(_01163_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06768_ (.I(_05824_),
    .Z(_01164_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06769_ (.A1(_01164_),
    .A2(_01011_),
    .B(_00556_),
    .ZN(_01165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _06770_ (.A1(_01161_),
    .A2(_00556_),
    .B1(_01163_),
    .B2(_01165_),
    .ZN(_01166_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06771_ (.A1(_01160_),
    .A2(_01166_),
    .Z(_01167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06772_ (.I(_01167_),
    .Z(_01168_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06773_ (.A1(_01099_),
    .A2(_00819_),
    .B(_01100_),
    .ZN(_01169_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06774_ (.A1(_01106_),
    .A2(_01113_),
    .Z(_01170_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06775_ (.A1(_01169_),
    .A2(_01170_),
    .ZN(_01171_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _06776_ (.A1(_01158_),
    .A2(_01168_),
    .A3(_01171_),
    .ZN(_01172_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06777_ (.I(_01160_),
    .Z(_01173_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06778_ (.A1(_01173_),
    .A2(_01166_),
    .Z(_01174_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06779_ (.A1(_01173_),
    .A2(_01166_),
    .ZN(_01175_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06780_ (.A1(_01174_),
    .A2(_01175_),
    .Z(_01176_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06781_ (.A1(_01158_),
    .A2(_01171_),
    .ZN(_01177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06782_ (.A1(_01176_),
    .A2(_01177_),
    .ZN(_01178_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06783_ (.A1(_01157_),
    .A2(_01172_),
    .A3(_01178_),
    .Z(_01179_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06784_ (.I(_00525_),
    .Z(_01180_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06785_ (.A1(_01180_),
    .A2(_00591_),
    .ZN(_01181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06786_ (.A1(_01181_),
    .A2(_01174_),
    .ZN(_01182_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06787_ (.A1(_01112_),
    .A2(_01175_),
    .B(_01182_),
    .C(_01121_),
    .ZN(_01183_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06788_ (.A1(_01068_),
    .A2(_01116_),
    .B(_01107_),
    .ZN(_01184_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06789_ (.A1(_01168_),
    .A2(_01184_),
    .Z(_01185_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06790_ (.A1(_01168_),
    .A2(_01184_),
    .B(_01126_),
    .ZN(_01186_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _06791_ (.A1(_01131_),
    .A2(_01176_),
    .B1(_01185_),
    .B2(_01186_),
    .ZN(_01187_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _06792_ (.A1(_01179_),
    .A2(_01183_),
    .A3(_01187_),
    .B1(_01173_),
    .B2(_01138_),
    .ZN(_01188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06793_ (.I(_01030_),
    .Z(_01189_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06794_ (.I(_01189_),
    .Z(_01190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06795_ (.I(_05827_),
    .Z(_01191_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06796_ (.A1(_01191_),
    .A2(_00443_),
    .Z(_01192_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06797_ (.I(\as2650.idx_ctrl[0] ),
    .ZN(_01193_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06798_ (.A1(_01009_),
    .A2(_01193_),
    .ZN(_01194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06799_ (.A1(_01009_),
    .A2(_01193_),
    .ZN(_01195_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06800_ (.A1(_05841_),
    .A2(_01194_),
    .B(_01195_),
    .ZN(_01196_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _06801_ (.A1(_01192_),
    .A2(_01196_),
    .Z(_01197_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06802_ (.A1(_01192_),
    .A2(_01196_),
    .ZN(_01198_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06803_ (.A1(_01197_),
    .A2(_01198_),
    .ZN(_01199_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _06804_ (.I(\as2650.addr_buff[5] ),
    .ZN(_01200_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06805_ (.A1(\as2650.addr_buff[6] ),
    .A2(_01200_),
    .ZN(_01201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06806_ (.A1(_01035_),
    .A2(_01200_),
    .ZN(_01202_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06807_ (.A1(_00443_),
    .A2(_01201_),
    .B(_01202_),
    .ZN(_01203_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06808_ (.A1(_01192_),
    .A2(_01203_),
    .Z(_01204_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06809_ (.A1(_01192_),
    .A2(_01203_),
    .ZN(_01205_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06810_ (.A1(_01204_),
    .A2(_01205_),
    .ZN(_01206_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06811_ (.A1(_01058_),
    .A2(_01206_),
    .ZN(_01207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06812_ (.I(_01164_),
    .Z(_01208_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06813_ (.I(_01208_),
    .Z(_01209_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06814_ (.A1(_00815_),
    .A2(_01021_),
    .A3(_01148_),
    .Z(_01210_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06815_ (.I(_05822_),
    .Z(_01211_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06816_ (.I(_01211_),
    .Z(_01212_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06817_ (.I(net9),
    .Z(_01213_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06818_ (.I(_01213_),
    .Z(_01214_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06819_ (.I(_01214_),
    .Z(_01215_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06820_ (.I(_01215_),
    .Z(_01216_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _06821_ (.A1(_00656_),
    .A2(_01000_),
    .A3(_01001_),
    .A4(_01004_),
    .ZN(_01217_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06822_ (.I(_01217_),
    .Z(_01218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06823_ (.A1(_00454_),
    .A2(_01218_),
    .ZN(_01219_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06824_ (.A1(_01216_),
    .A2(_01218_),
    .B(_01076_),
    .C(_01219_),
    .ZN(_01220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06825_ (.I(_01083_),
    .Z(_01221_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06826_ (.I(_01221_),
    .Z(_01222_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06827_ (.A1(_01212_),
    .A2(_01076_),
    .B(_01220_),
    .C(_01222_),
    .ZN(_01223_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06828_ (.I(_00445_),
    .Z(_01224_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06829_ (.I(_01224_),
    .Z(_01225_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06830_ (.A1(_01225_),
    .A2(_01064_),
    .B(_01210_),
    .ZN(_01226_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06831_ (.A1(_01209_),
    .A2(_01210_),
    .B1(_01223_),
    .B2(_01226_),
    .C(_01090_),
    .ZN(_01227_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06832_ (.A1(_01207_),
    .A2(_01227_),
    .B(_01097_),
    .ZN(_01228_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06833_ (.A1(_01190_),
    .A2(_01199_),
    .B(_01228_),
    .ZN(_01229_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06834_ (.I(_01008_),
    .Z(_01230_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06835_ (.I(_01018_),
    .Z(_01231_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _06836_ (.A1(_01230_),
    .A2(_01014_),
    .A3(_01015_),
    .A4(_01231_),
    .Z(_01232_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06837_ (.I0(net81),
    .I1(_01229_),
    .S(_01232_),
    .Z(_01233_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06838_ (.I(_01153_),
    .Z(_01234_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06839_ (.I0(\as2650.r123[0][1] ),
    .I1(\as2650.r123_2[0][1] ),
    .S(_05764_),
    .Z(_01235_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06840_ (.I(_01235_),
    .Z(_01236_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06841_ (.I(_01236_),
    .Z(_01237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06842_ (.A1(_01053_),
    .A2(_01237_),
    .ZN(_01238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06843_ (.A1(_01208_),
    .A2(_01145_),
    .ZN(_01239_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06844_ (.A1(_01238_),
    .A2(_01239_),
    .Z(_01240_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06845_ (.I(_01151_),
    .Z(_01241_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06846_ (.A1(\as2650.r123[1][1] ),
    .A2(_01234_),
    .B1(_01240_),
    .B2(_01241_),
    .ZN(_01242_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06847_ (.A1(_01156_),
    .A2(_01233_),
    .B(_01242_),
    .ZN(_00015_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06848_ (.I(_01194_),
    .Z(_01243_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06849_ (.I(_01195_),
    .Z(_01244_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _06850_ (.A1(_05821_),
    .A2(_01191_),
    .A3(_00443_),
    .Z(_01245_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _06851_ (.A1(_00431_),
    .A2(_00444_),
    .B(_00430_),
    .ZN(_01246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06852_ (.A1(_00430_),
    .A2(_01244_),
    .ZN(_01247_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _06853_ (.A1(_01244_),
    .A2(_01245_),
    .A3(_01246_),
    .B(_01247_),
    .ZN(_01248_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06854_ (.A1(_01243_),
    .A2(_01248_),
    .Z(_01249_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _06855_ (.A1(_05820_),
    .A2(_01191_),
    .A3(_05834_),
    .Z(_01250_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06856_ (.I(_01250_),
    .Z(_01251_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06857_ (.A1(_05828_),
    .A2(_00444_),
    .B(_05822_),
    .ZN(_01252_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06858_ (.A1(_01243_),
    .A2(_01251_),
    .A3(_01252_),
    .ZN(_01253_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _06859_ (.A1(_01249_),
    .A2(_01253_),
    .Z(_01254_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _06860_ (.A1(_01251_),
    .A2(_01252_),
    .B(_01035_),
    .C(_01200_),
    .ZN(_01255_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06861_ (.I(_01202_),
    .Z(_01256_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06862_ (.I(_01092_),
    .Z(_01257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06863_ (.A1(_00430_),
    .A2(_01257_),
    .ZN(_01258_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_4 _06864_ (.A1(_01256_),
    .A2(_01245_),
    .A3(_01246_),
    .B(_01258_),
    .ZN(_01259_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06865_ (.A1(_01255_),
    .A2(_01259_),
    .ZN(_01260_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06866_ (.I(_05850_),
    .Z(_01261_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06867_ (.I(_01261_),
    .Z(_01262_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06868_ (.I(_01074_),
    .Z(_01263_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _06869_ (.I(net10),
    .Z(_01264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06870_ (.I(_01264_),
    .Z(_01265_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06871_ (.I(_01217_),
    .Z(_01266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06872_ (.A1(_00450_),
    .A2(_01266_),
    .ZN(_01267_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06873_ (.A1(_01265_),
    .A2(_01218_),
    .B(_01077_),
    .C(_01267_),
    .ZN(_01268_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06874_ (.A1(_01262_),
    .A2(_01263_),
    .B(_01268_),
    .C(_01084_),
    .ZN(_01269_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06875_ (.A1(_01073_),
    .A2(_01222_),
    .B(_01269_),
    .ZN(_01270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06876_ (.I(_00438_),
    .Z(_01271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06877_ (.I(_01271_),
    .Z(_01272_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06878_ (.A1(_01272_),
    .A2(_01059_),
    .B(_01057_),
    .ZN(_01273_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06879_ (.A1(_01055_),
    .A2(_01270_),
    .B(_01273_),
    .ZN(_01274_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06880_ (.A1(_01090_),
    .A2(_01260_),
    .B(_01274_),
    .ZN(_01275_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06881_ (.I0(_01254_),
    .I1(_01275_),
    .S(_01097_),
    .Z(_01276_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _06882_ (.A1(_01110_),
    .A2(_00525_),
    .A3(_01118_),
    .ZN(_01277_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06883_ (.A1(_01158_),
    .A2(_01171_),
    .B(_01168_),
    .ZN(_01278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06884_ (.A1(\as2650.holding_reg[2] ),
    .A2(_00809_),
    .ZN(_01279_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06885_ (.A1(_01211_),
    .A2(_01105_),
    .B(_01279_),
    .ZN(_01280_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06886_ (.I(_01280_),
    .ZN(_01281_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06887_ (.I(_00440_),
    .ZN(_01282_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06888_ (.A1(_01282_),
    .A2(_01010_),
    .B1(_01011_),
    .B2(_01271_),
    .ZN(_01283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06889_ (.A1(\as2650.holding_reg[2] ),
    .A2(_00557_),
    .ZN(_01284_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06890_ (.A1(_00558_),
    .A2(_01283_),
    .B(_01284_),
    .ZN(_01285_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06891_ (.A1(_01281_),
    .A2(_01285_),
    .Z(_01286_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06892_ (.I(_01286_),
    .Z(_01287_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06893_ (.I(_01173_),
    .ZN(_01288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06894_ (.A1(_01288_),
    .A2(_01166_),
    .ZN(_01289_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06895_ (.I(_01289_),
    .ZN(_01290_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06896_ (.A1(_01278_),
    .A2(_01287_),
    .A3(_01290_),
    .ZN(_01291_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06897_ (.I(_01280_),
    .Z(_01292_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06898_ (.I(_01285_),
    .Z(_01293_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06899_ (.A1(_01292_),
    .A2(_01293_),
    .Z(_01294_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _06900_ (.A1(_01178_),
    .A2(_01289_),
    .B(_01294_),
    .ZN(_01295_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _06901_ (.A1(_01277_),
    .A2(_01291_),
    .A3(_01295_),
    .ZN(_01296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06902_ (.A1(_01292_),
    .A2(_01293_),
    .ZN(_01297_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06903_ (.A1(_01292_),
    .A2(_01293_),
    .ZN(_01298_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _06904_ (.A1(_01109_),
    .A2(_01297_),
    .B1(_01298_),
    .B2(_01112_),
    .C(_01121_),
    .ZN(_01299_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06905_ (.A1(_01167_),
    .A2(_01184_),
    .B(_01174_),
    .ZN(_01300_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06906_ (.A1(_01286_),
    .A2(_01300_),
    .Z(_01301_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06907_ (.A1(_01287_),
    .A2(_01300_),
    .B(_01127_),
    .ZN(_01302_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _06908_ (.A1(_01131_),
    .A2(_01287_),
    .B1(_01301_),
    .B2(_01302_),
    .ZN(_01303_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _06909_ (.A1(_01296_),
    .A2(_01299_),
    .A3(_01303_),
    .B1(_01292_),
    .B2(_01138_),
    .ZN(_01304_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06910_ (.I0(_01276_),
    .I1(net80),
    .S(_01019_),
    .Z(_01305_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06911_ (.A1(_01238_),
    .A2(_01239_),
    .Z(_01306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06912_ (.A1(_00438_),
    .A2(_01145_),
    .ZN(_01307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06913_ (.A1(_01164_),
    .A2(_01237_),
    .ZN(_01308_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06914_ (.A1(_01307_),
    .A2(_01308_),
    .ZN(_01309_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06915_ (.I0(\as2650.r123[0][2] ),
    .I1(\as2650.r123_2[0][2] ),
    .S(_05764_),
    .Z(_01310_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06916_ (.I(_01310_),
    .Z(_01311_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06917_ (.I(_01311_),
    .Z(_01312_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06918_ (.I(_01312_),
    .Z(_01313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06919_ (.A1(_01052_),
    .A2(_01313_),
    .ZN(_01314_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06920_ (.A1(_01309_),
    .A2(_01314_),
    .Z(_01315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06921_ (.A1(_01309_),
    .A2(_01314_),
    .ZN(_01316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06922_ (.A1(_01315_),
    .A2(_01316_),
    .ZN(_01317_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06923_ (.A1(_01306_),
    .A2(_01317_),
    .Z(_01318_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06924_ (.A1(\as2650.r123[1][2] ),
    .A2(_01234_),
    .B1(_01318_),
    .B2(_01241_),
    .ZN(_01319_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06925_ (.A1(_01156_),
    .A2(_01305_),
    .B(_01319_),
    .ZN(_00016_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06926_ (.A1(_05814_),
    .A2(_01250_),
    .Z(_01320_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _06927_ (.A1(_05849_),
    .A2(_01245_),
    .Z(_01321_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _06928_ (.A1(_01091_),
    .A2(_01036_),
    .ZN(_01322_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _06929_ (.A1(_05850_),
    .A2(_01257_),
    .B1(_01320_),
    .B2(_01201_),
    .C1(_01321_),
    .C2(_01322_),
    .ZN(_01323_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06930_ (.I(_05809_),
    .Z(_01324_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06931_ (.I(_01324_),
    .Z(_01325_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06932_ (.I(_01023_),
    .Z(_01326_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06933_ (.I(net11),
    .ZN(_01327_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06934_ (.I(_01327_),
    .Z(_01328_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06935_ (.A1(_00452_),
    .A2(_01005_),
    .Z(_01329_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06936_ (.A1(_01328_),
    .A2(_01218_),
    .B(_01075_),
    .C(_01329_),
    .ZN(_01330_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06937_ (.A1(_05805_),
    .A2(_01263_),
    .B(_01330_),
    .C(_01084_),
    .ZN(_01331_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _06938_ (.A1(_01211_),
    .A2(_01222_),
    .B(_01331_),
    .C(_01059_),
    .ZN(_01332_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06939_ (.A1(_01325_),
    .A2(_01326_),
    .B(_01332_),
    .ZN(_01333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06940_ (.A1(_01041_),
    .A2(_01333_),
    .ZN(_01334_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06941_ (.A1(_01041_),
    .A2(_01323_),
    .B(_01334_),
    .ZN(_01335_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06942_ (.I(_01189_),
    .Z(_01336_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06943_ (.I(_01244_),
    .Z(_01337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06944_ (.A1(_00434_),
    .A2(_01337_),
    .ZN(_01338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06945_ (.A1(_01048_),
    .A2(_01049_),
    .ZN(_01339_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06946_ (.I(_01339_),
    .Z(_01340_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _06947_ (.A1(_01337_),
    .A2(_01321_),
    .B(_01338_),
    .C(_01340_),
    .ZN(_01341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06948_ (.A1(_01243_),
    .A2(_01320_),
    .ZN(_01342_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _06949_ (.A1(_01341_),
    .A2(_01342_),
    .Z(_01343_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06950_ (.A1(_01336_),
    .A2(_01343_),
    .ZN(_01344_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _06951_ (.A1(_01190_),
    .A2(_01335_),
    .B(_01344_),
    .ZN(_01345_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06952_ (.I(_01120_),
    .Z(_01346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06953_ (.A1(\as2650.holding_reg[3] ),
    .A2(_00810_),
    .ZN(_01347_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06954_ (.A1(_01261_),
    .A2(_00810_),
    .B(_01347_),
    .ZN(_01348_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06955_ (.I(_01348_),
    .Z(_01349_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _06956_ (.I(_01110_),
    .Z(_01350_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06957_ (.I(_05813_),
    .ZN(_01351_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06958_ (.A1(_01351_),
    .A2(_01010_),
    .B1(_01011_),
    .B2(_01324_),
    .ZN(_01352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06959_ (.A1(\as2650.holding_reg[3] ),
    .A2(_00558_),
    .ZN(_01353_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06960_ (.A1(_00558_),
    .A2(_01352_),
    .B(_01353_),
    .ZN(_01354_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _06961_ (.A1(_01348_),
    .A2(_01354_),
    .Z(_01355_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06962_ (.I(_01354_),
    .Z(_01356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06963_ (.A1(_01349_),
    .A2(_01356_),
    .ZN(_01357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _06964_ (.A1(_01355_),
    .A2(_01357_),
    .ZN(_01358_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06965_ (.A1(_01286_),
    .A2(_01300_),
    .B(_01297_),
    .ZN(_01359_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06966_ (.A1(_01358_),
    .A2(_01359_),
    .Z(_01360_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _06967_ (.A1(_01350_),
    .A2(_01117_),
    .A3(_01360_),
    .ZN(_01361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06968_ (.I(_01277_),
    .Z(_01362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06969_ (.A1(_01281_),
    .A2(_01293_),
    .ZN(_01363_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06970_ (.I(_01363_),
    .ZN(_01364_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06971_ (.A1(_01295_),
    .A2(_01364_),
    .ZN(_01365_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _06972_ (.A1(_01358_),
    .A2(_01365_),
    .Z(_01366_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _06973_ (.A1(_01349_),
    .A2(_01356_),
    .Z(_01367_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _06974_ (.I(_01111_),
    .Z(_01368_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _06975_ (.A1(_01130_),
    .A2(_01367_),
    .B(_01368_),
    .ZN(_01369_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _06976_ (.A1(_00943_),
    .A2(_00961_),
    .A3(_01119_),
    .Z(_01370_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _06977_ (.A1(_01181_),
    .A2(_01367_),
    .B1(_01369_),
    .B2(_01355_),
    .C(_01370_),
    .ZN(_01371_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _06978_ (.A1(_01362_),
    .A2(_01366_),
    .B(_01371_),
    .ZN(_01372_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _06979_ (.A1(_01346_),
    .A2(_01349_),
    .B1(_01361_),
    .B2(_01372_),
    .ZN(_01373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06980_ (.A1(_01047_),
    .A2(_01373_),
    .ZN(_01374_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _06981_ (.A1(_01047_),
    .A2(_01345_),
    .B(_01374_),
    .ZN(_01375_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _06982_ (.A1(_01306_),
    .A2(_01317_),
    .ZN(_01376_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _06983_ (.A1(_01307_),
    .A2(_01308_),
    .Z(_01377_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _06984_ (.I(_01377_),
    .ZN(_01378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06985_ (.A1(_05807_),
    .A2(_01145_),
    .ZN(_01379_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _06986_ (.I(_05815_),
    .Z(_01380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _06987_ (.A1(_01380_),
    .A2(_01236_),
    .ZN(_01381_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _06988_ (.A1(_01379_),
    .A2(_01381_),
    .ZN(_01382_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06989_ (.I(\as2650.r0[1] ),
    .Z(_01383_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _06990_ (.I0(\as2650.r123[0][3] ),
    .I1(\as2650.r123_2[0][3] ),
    .S(net51),
    .Z(_01384_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06991_ (.I(_01384_),
    .Z(_01385_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06992_ (.I(_01310_),
    .Z(_01386_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _06993_ (.A1(_01383_),
    .A2(\as2650.r0[0] ),
    .A3(_01385_),
    .A4(_01386_),
    .Z(_01387_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06994_ (.I(_01387_),
    .Z(_01388_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _06995_ (.I(_01384_),
    .Z(_01389_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _06996_ (.I(_01389_),
    .Z(_01390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _06997_ (.I(_01390_),
    .Z(_01391_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _06998_ (.A1(_05830_),
    .A2(_01391_),
    .B1(_01313_),
    .B2(_05824_),
    .ZN(_01392_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _06999_ (.A1(_01388_),
    .A2(_01392_),
    .ZN(_01393_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07000_ (.A1(_01382_),
    .A2(_01393_),
    .Z(_01394_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07001_ (.A1(_01315_),
    .A2(_01394_),
    .Z(_01395_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07002_ (.A1(_01377_),
    .A2(_01394_),
    .Z(_01396_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07003_ (.A1(_01378_),
    .A2(_01395_),
    .B(_01396_),
    .ZN(_01397_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07004_ (.A1(_01376_),
    .A2(_01397_),
    .Z(_01398_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _07005_ (.A1(_05744_),
    .A2(_00566_),
    .A3(_00821_),
    .ZN(_01399_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07006_ (.I(_01148_),
    .Z(_01400_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07007_ (.A1(_01147_),
    .A2(_01399_),
    .A3(_01400_),
    .ZN(_01401_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07008_ (.I(_01401_),
    .Z(_01402_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07009_ (.I(_01402_),
    .Z(_01403_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07010_ (.A1(\as2650.r123[1][3] ),
    .A2(_01154_),
    .ZN(_01404_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07011_ (.A1(_01046_),
    .A2(_01375_),
    .B1(_01398_),
    .B2(_01403_),
    .C(_01404_),
    .ZN(_00017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07012_ (.I(_01339_),
    .Z(_01405_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07013_ (.A1(_05849_),
    .A2(_01250_),
    .ZN(_01406_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _07014_ (.A1(_05847_),
    .A2(_01406_),
    .Z(_01407_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _07015_ (.A1(_05849_),
    .A2(_05821_),
    .A3(_01191_),
    .A4(_05834_),
    .ZN(_01408_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07016_ (.A1(_05847_),
    .A2(_01408_),
    .Z(_01409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07017_ (.A1(_05848_),
    .A2(_01244_),
    .ZN(_01410_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07018_ (.A1(_01337_),
    .A2(_01409_),
    .B(_01410_),
    .C(_01405_),
    .ZN(_01411_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07019_ (.A1(_01405_),
    .A2(_01407_),
    .B(_01411_),
    .ZN(_01412_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07020_ (.I(_01412_),
    .Z(_01413_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07021_ (.A1(_01256_),
    .A2(_01409_),
    .ZN(_01414_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _07022_ (.A1(_05848_),
    .A2(_01257_),
    .B1(_01407_),
    .B2(_01201_),
    .C(_01414_),
    .ZN(_01415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07023_ (.I(_01415_),
    .Z(_01416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07024_ (.A1(_01090_),
    .A2(_01416_),
    .ZN(_01417_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07025_ (.I(_05797_),
    .Z(_01418_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07026_ (.I(_01418_),
    .Z(_01419_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07027_ (.I(_01419_),
    .Z(_01420_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07028_ (.I(_01420_),
    .Z(_01421_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07029_ (.I(_00425_),
    .Z(_01422_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07030_ (.I(net12),
    .Z(_01423_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07031_ (.I(_01423_),
    .Z(_01424_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07032_ (.I(_01424_),
    .Z(_01425_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07033_ (.I(_01425_),
    .Z(_01426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07034_ (.A1(_01426_),
    .A2(_01006_),
    .ZN(_01427_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07035_ (.A1(_00437_),
    .A2(_01006_),
    .B(_01077_),
    .C(_01427_),
    .ZN(_01428_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07036_ (.I(_01221_),
    .Z(_01429_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07037_ (.A1(_01422_),
    .A2(_01076_),
    .B(_01428_),
    .C(_01429_),
    .ZN(_01430_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07038_ (.A1(_01262_),
    .A2(_01222_),
    .B(_01430_),
    .C(_01326_),
    .ZN(_01431_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07039_ (.A1(_01421_),
    .A2(_01055_),
    .B(_01058_),
    .C(_01431_),
    .ZN(_01432_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07040_ (.A1(_01336_),
    .A2(_01417_),
    .A3(_01432_),
    .ZN(_01433_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07041_ (.A1(_01190_),
    .A2(_01413_),
    .B(_01433_),
    .ZN(_01434_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07042_ (.A1(\as2650.holding_reg[4] ),
    .A2(_00810_),
    .ZN(_01435_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _07043_ (.A1(_00429_),
    .A2(_00811_),
    .B(_01435_),
    .ZN(_01436_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07044_ (.I(_05803_),
    .ZN(_01437_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _07045_ (.A1(_01437_),
    .A2(_01025_),
    .B1(_01012_),
    .B2(_01419_),
    .ZN(_01438_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07046_ (.A1(\as2650.holding_reg[4] ),
    .A2(_00819_),
    .ZN(_01439_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _07047_ (.A1(_00819_),
    .A2(_01438_),
    .B(_01439_),
    .ZN(_01440_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07048_ (.A1(_01436_),
    .A2(_01440_),
    .ZN(_01441_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07049_ (.I(_01441_),
    .ZN(_01442_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07050_ (.A1(_01436_),
    .A2(_01440_),
    .ZN(_01443_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07051_ (.A1(_01442_),
    .A2(_01443_),
    .ZN(_01444_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07052_ (.A1(_01355_),
    .A2(_01359_),
    .B(_01367_),
    .ZN(_01445_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07053_ (.A1(_01444_),
    .A2(_01445_),
    .Z(_01446_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07054_ (.A1(_01127_),
    .A2(_01446_),
    .Z(_01447_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07055_ (.A1(_01278_),
    .A2(_01290_),
    .B(_01286_),
    .ZN(_01448_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _07056_ (.A1(_01355_),
    .A2(_01357_),
    .B1(_01363_),
    .B2(_01448_),
    .ZN(_01449_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07057_ (.I(_01349_),
    .ZN(_01450_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07058_ (.A1(_01450_),
    .A2(_01356_),
    .Z(_01451_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07059_ (.A1(_01449_),
    .A2(_01444_),
    .A3(_01451_),
    .ZN(_01452_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07060_ (.A1(_01449_),
    .A2(_01451_),
    .B(_01444_),
    .ZN(_01453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07061_ (.A1(_01157_),
    .A2(_01453_),
    .ZN(_01454_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07062_ (.A1(_01452_),
    .A2(_01454_),
    .ZN(_01455_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07063_ (.I(_01370_),
    .Z(_01456_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _07064_ (.A1(_01368_),
    .A2(_01441_),
    .B1(_01443_),
    .B2(_01109_),
    .ZN(_01457_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07065_ (.A1(_01456_),
    .A2(_01457_),
    .ZN(_01458_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07066_ (.A1(_01131_),
    .A2(_01444_),
    .B(_01458_),
    .ZN(_01459_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _07067_ (.A1(_01447_),
    .A2(_01455_),
    .A3(_01459_),
    .B1(_01436_),
    .B2(_01346_),
    .ZN(_01460_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07068_ (.I(_01460_),
    .Z(_01461_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07069_ (.I0(_01434_),
    .I1(_01461_),
    .S(_01019_),
    .Z(_01462_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07070_ (.I(_01397_),
    .ZN(_01463_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07071_ (.A1(_01376_),
    .A2(_01463_),
    .ZN(_01464_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07072_ (.A1(_01377_),
    .A2(_01315_),
    .B(_01394_),
    .ZN(_01465_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07073_ (.A1(_01379_),
    .A2(_01381_),
    .Z(_01466_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07074_ (.I0(\as2650.r123[0][4] ),
    .I1(\as2650.r123_2[0][4] ),
    .S(_05799_),
    .Z(_01467_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07075_ (.I(_01467_),
    .Z(_01468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07076_ (.A1(_01052_),
    .A2(_01468_),
    .ZN(_01469_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07077_ (.A1(_01466_),
    .A2(_01469_),
    .Z(_01470_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _07078_ (.A1(_01382_),
    .A2(_01388_),
    .A3(_01392_),
    .Z(_01471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07079_ (.I(_01235_),
    .Z(_01472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07080_ (.A1(\as2650.r0[3] ),
    .A2(_01472_),
    .ZN(_01473_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07081_ (.A1(\as2650.r0[4] ),
    .A2(_01144_),
    .ZN(_01474_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07082_ (.A1(_01473_),
    .A2(_01474_),
    .Z(_01475_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07083_ (.I(_01390_),
    .Z(_01476_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _07084_ (.A1(_05824_),
    .A2(_01476_),
    .B1(_01312_),
    .B2(_01380_),
    .ZN(_01477_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07085_ (.I(_01477_),
    .ZN(_01478_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _07086_ (.A1(_01380_),
    .A2(_05823_),
    .A3(_01476_),
    .A4(_01312_),
    .ZN(_01479_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07087_ (.A1(_01388_),
    .A2(_01479_),
    .Z(_01480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07088_ (.A1(_01478_),
    .A2(_01480_),
    .ZN(_01481_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07089_ (.A1(_01471_),
    .A2(_01475_),
    .A3(_01481_),
    .Z(_01482_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07090_ (.A1(_01470_),
    .A2(_01482_),
    .Z(_01483_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07091_ (.A1(_01465_),
    .A2(_01483_),
    .Z(_01484_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07092_ (.A1(_01464_),
    .A2(_01484_),
    .Z(_01485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07093_ (.A1(\as2650.r123[1][4] ),
    .A2(_01154_),
    .ZN(_01486_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07094_ (.A1(_01046_),
    .A2(_01462_),
    .B1(_01485_),
    .B2(_01403_),
    .C(_01486_),
    .ZN(_00018_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07095_ (.I(_01232_),
    .Z(_01487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07096_ (.A1(_00425_),
    .A2(_00559_),
    .ZN(_01488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07097_ (.A1(\as2650.holding_reg[5] ),
    .A2(_00811_),
    .ZN(_01489_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07098_ (.A1(_01488_),
    .A2(_01489_),
    .Z(_01490_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07099_ (.A1(_01488_),
    .A2(_01489_),
    .ZN(_01491_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07100_ (.I(_05794_),
    .ZN(_01492_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07101_ (.I(_05787_),
    .Z(_01493_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _07102_ (.A1(_01492_),
    .A2(_01025_),
    .B1(_01012_),
    .B2(_01493_),
    .ZN(_01494_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07103_ (.A1(\as2650.holding_reg[5] ),
    .A2(_00559_),
    .ZN(_01495_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07104_ (.A1(_00559_),
    .A2(_01494_),
    .B(_01495_),
    .ZN(_01496_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07105_ (.A1(_01491_),
    .A2(_01496_),
    .Z(_01497_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07106_ (.I(_01497_),
    .Z(_01498_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07107_ (.I(_00429_),
    .Z(_01499_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _07108_ (.A1(_01499_),
    .A2(_00812_),
    .B(_01435_),
    .C(_01440_),
    .ZN(_01500_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07109_ (.A1(_01453_),
    .A2(_01498_),
    .A3(_01500_),
    .ZN(_01501_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07110_ (.A1(_01453_),
    .A2(_01500_),
    .B(_01497_),
    .ZN(_01502_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07111_ (.A1(_01362_),
    .A2(_01502_),
    .ZN(_01503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07112_ (.A1(_01501_),
    .A2(_01503_),
    .ZN(_01504_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07113_ (.I(_01127_),
    .Z(_01505_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07114_ (.A1(_01443_),
    .A2(_01445_),
    .B(_01441_),
    .ZN(_01506_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07115_ (.A1(_01498_),
    .A2(_01506_),
    .Z(_01507_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07116_ (.A1(_01491_),
    .A2(_01496_),
    .Z(_01508_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07117_ (.A1(_01491_),
    .A2(_01496_),
    .Z(_01509_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07118_ (.A1(_01130_),
    .A2(_01508_),
    .B(_01112_),
    .ZN(_01510_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07119_ (.A1(_01181_),
    .A2(_01508_),
    .B1(_01509_),
    .B2(_01510_),
    .ZN(_01511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07120_ (.A1(_01346_),
    .A2(_01511_),
    .ZN(_01512_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07121_ (.A1(_01505_),
    .A2(_01507_),
    .B(_01512_),
    .ZN(_01513_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _07122_ (.A1(_01456_),
    .A2(_01490_),
    .B1(_01504_),
    .B2(_01513_),
    .ZN(_01514_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07123_ (.I(_01340_),
    .Z(_01515_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07124_ (.A1(_05840_),
    .A2(_05804_),
    .A3(_01406_),
    .ZN(_01516_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _07125_ (.A1(_00429_),
    .A2(_01261_),
    .A3(_01251_),
    .B(_05795_),
    .ZN(_01517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07126_ (.A1(_01516_),
    .A2(_01517_),
    .ZN(_01518_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07127_ (.I(_01337_),
    .Z(_01519_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07128_ (.A1(_05805_),
    .A2(_01408_),
    .ZN(_01520_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07129_ (.A1(_05840_),
    .A2(_01520_),
    .Z(_01521_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07130_ (.I(_05795_),
    .Z(_01522_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07131_ (.A1(_01522_),
    .A2(_01519_),
    .ZN(_01523_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07132_ (.A1(_01519_),
    .A2(_01521_),
    .B(_01523_),
    .C(_01515_),
    .ZN(_01524_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07133_ (.A1(_01515_),
    .A2(_01518_),
    .B(_01524_),
    .ZN(_01525_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07134_ (.I(_01525_),
    .Z(_01526_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07135_ (.I(_01257_),
    .Z(_01527_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07136_ (.I(_01201_),
    .Z(_01528_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07137_ (.A1(_01256_),
    .A2(_01521_),
    .ZN(_01529_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _07138_ (.A1(_01522_),
    .A2(_01527_),
    .B1(_01518_),
    .B2(_01528_),
    .C(_01529_),
    .ZN(_01530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07139_ (.I(_01530_),
    .Z(_01531_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07140_ (.A1(_01089_),
    .A2(_01531_),
    .ZN(_01532_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07141_ (.I(_01493_),
    .Z(_01533_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07142_ (.I(_00422_),
    .Z(_01534_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _07143_ (.I(net1),
    .ZN(_01535_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07144_ (.I(_01535_),
    .Z(_01536_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07145_ (.A1(_00428_),
    .A2(_01217_),
    .ZN(_01537_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07146_ (.A1(_01536_),
    .A2(_01266_),
    .B(_01075_),
    .C(_01537_),
    .ZN(_01538_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07147_ (.A1(_01534_),
    .A2(_01263_),
    .B(_01538_),
    .C(_01084_),
    .ZN(_01539_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07148_ (.A1(_01499_),
    .A2(_01429_),
    .B(_01539_),
    .C(_01059_),
    .ZN(_01540_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07149_ (.A1(_01533_),
    .A2(_01055_),
    .B(_01058_),
    .C(_01540_),
    .ZN(_01541_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07150_ (.A1(_01097_),
    .A2(_01532_),
    .A3(_01541_),
    .ZN(_01542_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07151_ (.A1(_01190_),
    .A2(_01526_),
    .B(_01542_),
    .ZN(_01543_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07152_ (.A1(_01487_),
    .A2(_01543_),
    .ZN(_01544_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _07153_ (.A1(_01487_),
    .A2(_01514_),
    .B(_01544_),
    .ZN(_01545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07154_ (.A1(_01465_),
    .A2(_01483_),
    .ZN(_01546_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07155_ (.A1(_01376_),
    .A2(_01463_),
    .A3(_01484_),
    .ZN(_01547_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07156_ (.A1(_01466_),
    .A2(_01469_),
    .ZN(_01548_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07157_ (.A1(_01473_),
    .A2(_01474_),
    .ZN(_01549_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07158_ (.A1(_01549_),
    .A2(_01478_),
    .A3(_01480_),
    .ZN(_01550_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _07159_ (.A1(_05816_),
    .A2(_05823_),
    .A3(_01385_),
    .A4(_01386_),
    .Z(_01551_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07160_ (.A1(_01387_),
    .A2(_01551_),
    .Z(_01552_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07161_ (.A1(_01477_),
    .A2(_01552_),
    .B(_01475_),
    .ZN(_01553_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07162_ (.A1(_01550_),
    .A2(_01553_),
    .B(_01471_),
    .ZN(_01554_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07163_ (.A1(_01470_),
    .A2(_01482_),
    .B(_01554_),
    .ZN(_01555_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07164_ (.A1(_01473_),
    .A2(_01474_),
    .ZN(_01556_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07165_ (.I0(\as2650.r123[0][5] ),
    .I1(\as2650.r123_2[0][5] ),
    .S(_05774_),
    .Z(_01557_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07166_ (.A1(_05830_),
    .A2(_01557_),
    .ZN(_01558_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07167_ (.A1(_01556_),
    .A2(_01558_),
    .ZN(_01559_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07168_ (.A1(_01164_),
    .A2(_01468_),
    .ZN(_01560_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07169_ (.A1(_01559_),
    .A2(_01560_),
    .Z(_01561_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07170_ (.A1(_01388_),
    .A2(_01479_),
    .ZN(_01562_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _07171_ (.A1(_01549_),
    .A2(_01477_),
    .A3(_01552_),
    .B(_01562_),
    .ZN(_01563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07172_ (.A1(\as2650.r0[4] ),
    .A2(_01472_),
    .ZN(_01564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07173_ (.A1(_05786_),
    .A2(_01143_),
    .ZN(_01565_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07174_ (.A1(_01564_),
    .A2(_01565_),
    .ZN(_01566_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _07175_ (.A1(\as2650.r0[3] ),
    .A2(_05815_),
    .A3(_01385_),
    .A4(_01310_),
    .ZN(_01567_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07176_ (.I(_01567_),
    .Z(_01568_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07177_ (.A1(_01551_),
    .A2(_01568_),
    .ZN(_01569_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _07178_ (.A1(_01380_),
    .A2(_01476_),
    .B1(_01311_),
    .B2(_05806_),
    .ZN(_01570_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07179_ (.A1(_01551_),
    .A2(_01568_),
    .Z(_01571_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07180_ (.A1(_01569_),
    .A2(_01570_),
    .A3(_01571_),
    .ZN(_01572_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07181_ (.A1(_01563_),
    .A2(_01566_),
    .A3(_01572_),
    .Z(_01573_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07182_ (.A1(_01561_),
    .A2(_01573_),
    .ZN(_01574_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _07183_ (.A1(_01548_),
    .A2(_01555_),
    .A3(_01574_),
    .ZN(_01575_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07184_ (.A1(_01546_),
    .A2(_01547_),
    .B(_01575_),
    .ZN(_01576_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07185_ (.A1(_01546_),
    .A2(_01547_),
    .A3(_01575_),
    .Z(_01577_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07186_ (.A1(_01576_),
    .A2(_01577_),
    .ZN(_01578_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07187_ (.A1(\as2650.r123[1][5] ),
    .A2(_01234_),
    .B1(_01578_),
    .B2(_01241_),
    .ZN(_01579_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07188_ (.A1(_01156_),
    .A2(_01545_),
    .B(_01579_),
    .ZN(_00019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07189_ (.I(_05861_),
    .Z(_01580_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07190_ (.I(_01580_),
    .Z(_01581_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07191_ (.I(_00811_),
    .Z(_01582_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07192_ (.A1(\as2650.holding_reg[6] ),
    .A2(_01582_),
    .ZN(_01583_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07193_ (.A1(_01581_),
    .A2(_01582_),
    .B(_01583_),
    .ZN(_01584_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07194_ (.I(_01584_),
    .ZN(_01585_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07195_ (.I(_05860_),
    .ZN(_01586_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07196_ (.I(_05855_),
    .Z(_01587_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _07197_ (.A1(_01586_),
    .A2(_01025_),
    .B1(_01012_),
    .B2(_01587_),
    .ZN(_01588_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07198_ (.A1(\as2650.holding_reg[6] ),
    .A2(_00820_),
    .ZN(_01589_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07199_ (.A1(_00820_),
    .A2(_01588_),
    .B(_01589_),
    .ZN(_01590_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _07200_ (.A1(_01584_),
    .A2(_01590_),
    .Z(_01591_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07201_ (.A1(_01584_),
    .A2(_01590_),
    .ZN(_01592_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07202_ (.A1(_01591_),
    .A2(_01592_),
    .ZN(_01593_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07203_ (.I(_01593_),
    .Z(_01594_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07204_ (.A1(_01490_),
    .A2(_01496_),
    .Z(_01595_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _07205_ (.A1(_01502_),
    .A2(_01594_),
    .A3(_01595_),
    .Z(_01596_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07206_ (.A1(_01502_),
    .A2(_01595_),
    .B(_01593_),
    .ZN(_01597_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07207_ (.A1(_01157_),
    .A2(_01596_),
    .A3(_01597_),
    .ZN(_01598_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07208_ (.A1(_01508_),
    .A2(_01506_),
    .B(_01509_),
    .ZN(_01599_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07209_ (.A1(_01594_),
    .A2(_01599_),
    .Z(_01600_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07210_ (.I(_00997_),
    .Z(_01601_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07211_ (.A1(_01601_),
    .A2(_01592_),
    .B(_01350_),
    .C(_00589_),
    .ZN(_01602_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07212_ (.I(_01591_),
    .ZN(_01603_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _07213_ (.A1(_01109_),
    .A2(_01592_),
    .B1(_01602_),
    .B2(_01603_),
    .C(_01138_),
    .ZN(_01604_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07214_ (.A1(_01505_),
    .A2(_01600_),
    .B(_01604_),
    .ZN(_01605_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _07215_ (.A1(_01456_),
    .A2(_01585_),
    .B1(_01598_),
    .B2(_01605_),
    .ZN(_01606_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _07216_ (.A1(_00422_),
    .A2(_01516_),
    .Z(_01607_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07217_ (.A1(_01048_),
    .A2(_01049_),
    .ZN(_01608_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _07218_ (.A1(_05839_),
    .A2(_05804_),
    .A3(_01408_),
    .ZN(_01609_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _07219_ (.A1(_05861_),
    .A2(_01609_),
    .Z(_01610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07220_ (.A1(_01608_),
    .A2(_01610_),
    .ZN(_01611_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07221_ (.A1(_00422_),
    .A2(_01608_),
    .B(_01611_),
    .C(_01340_),
    .ZN(_01612_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _07222_ (.A1(_01340_),
    .A2(_01607_),
    .B(_01612_),
    .ZN(_01613_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07223_ (.I(_01613_),
    .Z(_01614_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07224_ (.I(_01587_),
    .Z(_01615_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07225_ (.I(_01615_),
    .Z(_01616_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07226_ (.I(_01522_),
    .Z(_01617_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07227_ (.A1(_05768_),
    .A2(_05779_),
    .A3(_05784_),
    .ZN(_01618_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07228_ (.A1(_00424_),
    .A2(_01266_),
    .ZN(_01619_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07229_ (.I(net2),
    .Z(_01620_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07230_ (.I(_01620_),
    .Z(_01621_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07231_ (.I(_01621_),
    .Z(_01622_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07232_ (.I(_01622_),
    .Z(_01623_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07233_ (.I(_01623_),
    .Z(_01624_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07234_ (.A1(_01624_),
    .A2(_01005_),
    .ZN(_01625_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07235_ (.A1(_01075_),
    .A2(_01619_),
    .A3(_01625_),
    .ZN(_01626_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07236_ (.A1(_01618_),
    .A2(_01263_),
    .B(_01626_),
    .C(_01221_),
    .ZN(_01627_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07237_ (.A1(_01617_),
    .A2(_01429_),
    .B(_01627_),
    .C(_01024_),
    .ZN(_01628_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07238_ (.A1(_01616_),
    .A2(_01326_),
    .B(_01057_),
    .C(_01628_),
    .ZN(_01629_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _07239_ (.A1(_01580_),
    .A2(_01527_),
    .B1(_01607_),
    .B2(_01528_),
    .C1(_01610_),
    .C2(_01322_),
    .ZN(_01630_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07240_ (.I(_01630_),
    .Z(_01631_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07241_ (.A1(_01089_),
    .A2(_01631_),
    .ZN(_01632_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07242_ (.A1(_01189_),
    .A2(_01629_),
    .A3(_01632_),
    .ZN(_01633_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07243_ (.A1(_01336_),
    .A2(_01614_),
    .B(_01633_),
    .ZN(_01634_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07244_ (.A1(_01232_),
    .A2(_01634_),
    .ZN(_01635_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _07245_ (.A1(_01487_),
    .A2(_01606_),
    .B(_01635_),
    .ZN(_01636_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07246_ (.A1(_01555_),
    .A2(_01574_),
    .ZN(_01637_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07247_ (.A1(_01555_),
    .A2(_01574_),
    .ZN(_01638_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07248_ (.A1(_01548_),
    .A2(_01637_),
    .B(_01638_),
    .ZN(_01639_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07249_ (.I(_01468_),
    .Z(_01640_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07250_ (.A1(_01208_),
    .A2(_01640_),
    .A3(_01559_),
    .ZN(_01641_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _07251_ (.A1(_01473_),
    .A2(_01474_),
    .A3(_01558_),
    .B(_01641_),
    .ZN(_01642_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _07252_ (.A1(_01566_),
    .A2(_01569_),
    .A3(_01570_),
    .A4(_01571_),
    .Z(_01643_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _07253_ (.A1(_01569_),
    .A2(_01570_),
    .A3(_01571_),
    .B(_01566_),
    .ZN(_01644_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07254_ (.A1(_01563_),
    .A2(_01643_),
    .A3(_01644_),
    .ZN(_01645_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07255_ (.A1(_01561_),
    .A2(_01573_),
    .B(_01645_),
    .ZN(_01646_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07256_ (.A1(_01564_),
    .A2(_01565_),
    .ZN(_01647_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07257_ (.A1(_05823_),
    .A2(_01557_),
    .ZN(_01648_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07258_ (.A1(_01647_),
    .A2(_01648_),
    .ZN(_01649_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07259_ (.A1(_05817_),
    .A2(_01467_),
    .ZN(_01650_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07260_ (.A1(_01649_),
    .A2(_01650_),
    .Z(_01651_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07261_ (.A1(_01551_),
    .A2(_01568_),
    .ZN(_01652_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _07262_ (.A1(_01566_),
    .A2(_01569_),
    .A3(_01570_),
    .B(_01652_),
    .ZN(_01653_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07263_ (.I0(\as2650.r123[0][6] ),
    .I1(\as2650.r123_2[0][6] ),
    .S(_05764_),
    .Z(_01654_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07264_ (.A1(\as2650.r0[0] ),
    .A2(_01654_),
    .Z(_01655_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07265_ (.A1(\as2650.r0[5] ),
    .A2(_01472_),
    .ZN(_01656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07266_ (.A1(_05854_),
    .A2(_01144_),
    .ZN(_01657_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _07267_ (.A1(_01655_),
    .A2(_01656_),
    .A3(_01657_),
    .ZN(_01658_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _07268_ (.A1(_05807_),
    .A2(_01391_),
    .B1(_01312_),
    .B2(_05796_),
    .ZN(_01659_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _07269_ (.A1(_05796_),
    .A2(_05806_),
    .A3(_01390_),
    .A4(_01311_),
    .ZN(_01660_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07270_ (.A1(_01567_),
    .A2(_01660_),
    .Z(_01661_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07271_ (.A1(_01659_),
    .A2(_01661_),
    .ZN(_01662_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07272_ (.A1(_01653_),
    .A2(_01658_),
    .A3(_01662_),
    .Z(_01663_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07273_ (.A1(_01651_),
    .A2(_01663_),
    .Z(_01664_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07274_ (.A1(_01646_),
    .A2(_01664_),
    .Z(_01665_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07275_ (.A1(_01642_),
    .A2(_01665_),
    .ZN(_01666_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07276_ (.A1(_01639_),
    .A2(_01666_),
    .Z(_01667_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07277_ (.A1(_01576_),
    .A2(_01667_),
    .Z(_01668_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07278_ (.A1(\as2650.r123[1][6] ),
    .A2(_01234_),
    .B1(_01668_),
    .B2(_01241_),
    .ZN(_01669_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07279_ (.A1(_01156_),
    .A2(_01636_),
    .B(_01669_),
    .ZN(_00020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07280_ (.A1(\as2650.holding_reg[7] ),
    .A2(_01582_),
    .ZN(_01670_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07281_ (.A1(_01066_),
    .A2(_01582_),
    .B(_01670_),
    .ZN(_01671_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _07282_ (.I(_01671_),
    .ZN(_01672_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07283_ (.I(_05758_),
    .Z(_01673_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07284_ (.I(_01673_),
    .Z(_01674_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07285_ (.A1(_01066_),
    .A2(_01026_),
    .ZN(_01675_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _07286_ (.A1(_01674_),
    .A2(_01026_),
    .B(_01675_),
    .C(_00812_),
    .ZN(_01676_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07287_ (.A1(\as2650.holding_reg[7] ),
    .A2(_00560_),
    .ZN(_01677_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07288_ (.A1(_01676_),
    .A2(_01677_),
    .B(_01672_),
    .ZN(_01678_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07289_ (.I(_01678_),
    .ZN(_01679_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07290_ (.A1(_01672_),
    .A2(_01676_),
    .A3(_01677_),
    .ZN(_01680_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07291_ (.A1(_01679_),
    .A2(_01680_),
    .Z(_01681_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07292_ (.A1(_01585_),
    .A2(_01590_),
    .ZN(_01682_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _07293_ (.A1(_01597_),
    .A2(_01681_),
    .A3(_01682_),
    .Z(_01683_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07294_ (.A1(_01597_),
    .A2(_01682_),
    .B(_01681_),
    .ZN(_01684_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _07295_ (.A1(_01362_),
    .A2(_01683_),
    .A3(_01684_),
    .Z(_01685_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07296_ (.A1(_01592_),
    .A2(_01599_),
    .B(_01603_),
    .ZN(_01686_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07297_ (.A1(_01681_),
    .A2(_01686_),
    .Z(_01687_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07298_ (.I(_01678_),
    .Z(_01688_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07299_ (.I(_01680_),
    .Z(_01689_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07300_ (.A1(_01130_),
    .A2(_01688_),
    .B(_01368_),
    .ZN(_01690_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07301_ (.A1(_01181_),
    .A2(_01688_),
    .B1(_01689_),
    .B2(_01690_),
    .ZN(_01691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07302_ (.A1(_01121_),
    .A2(_01691_),
    .ZN(_01692_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07303_ (.A1(_01505_),
    .A2(_01687_),
    .B(_01692_),
    .ZN(_01693_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _07304_ (.A1(_01456_),
    .A2(_01672_),
    .B1(_01685_),
    .B2(_01693_),
    .ZN(_01694_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07305_ (.A1(_01580_),
    .A2(_01516_),
    .ZN(_01695_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _07306_ (.A1(_05785_),
    .A2(_01695_),
    .Z(_01696_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07307_ (.A1(_01580_),
    .A2(_01609_),
    .Z(_01697_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07308_ (.A1(_01618_),
    .A2(_01697_),
    .Z(_01698_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07309_ (.A1(_01066_),
    .A2(_01519_),
    .ZN(_01699_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07310_ (.A1(_01519_),
    .A2(_01698_),
    .B(_01699_),
    .C(_01515_),
    .ZN(_01700_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _07311_ (.A1(_01515_),
    .A2(_01696_),
    .B(_01700_),
    .ZN(_01701_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07312_ (.I(_01701_),
    .Z(_01702_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07313_ (.I(_01674_),
    .Z(_01703_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07314_ (.A1(_01065_),
    .A2(_01224_),
    .B(_01069_),
    .ZN(_01704_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_4 _07315_ (.I(_00847_),
    .ZN(_01705_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07316_ (.A1(_00421_),
    .A2(_01217_),
    .ZN(_01706_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _07317_ (.A1(_01705_),
    .A2(_01266_),
    .B(_01074_),
    .C(_01706_),
    .ZN(_01707_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07318_ (.A1(_01077_),
    .A2(_01704_),
    .B(_01707_),
    .C(_01221_),
    .ZN(_01708_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07319_ (.A1(_01581_),
    .A2(_01429_),
    .B(_01708_),
    .C(_01024_),
    .ZN(_01709_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _07320_ (.A1(_01703_),
    .A2(_01326_),
    .B(_01057_),
    .C(_01709_),
    .ZN(_01710_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07321_ (.A1(_01256_),
    .A2(_01698_),
    .ZN(_01711_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _07322_ (.A1(_01067_),
    .A2(_01527_),
    .B1(_01696_),
    .B2(_01528_),
    .C(_01711_),
    .ZN(_01712_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07323_ (.I(_01712_),
    .Z(_01713_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07324_ (.A1(_01089_),
    .A2(_01713_),
    .ZN(_01714_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07325_ (.A1(_01189_),
    .A2(_01710_),
    .A3(_01714_),
    .ZN(_01715_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07326_ (.A1(_01336_),
    .A2(_01702_),
    .B(_01715_),
    .ZN(_01716_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07327_ (.A1(_01232_),
    .A2(_01716_),
    .ZN(_01717_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _07328_ (.A1(_01487_),
    .A2(_01694_),
    .B(_01717_),
    .ZN(_01718_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07329_ (.A1(_01639_),
    .A2(_01666_),
    .ZN(_01719_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07330_ (.A1(_01576_),
    .A2(_01667_),
    .B(_01719_),
    .ZN(_01720_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07331_ (.A1(_01646_),
    .A2(_01664_),
    .ZN(_01721_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07332_ (.A1(_01642_),
    .A2(_01665_),
    .ZN(_01722_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07333_ (.A1(_01721_),
    .A2(_01722_),
    .ZN(_01723_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07334_ (.I(_01640_),
    .Z(_01724_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07335_ (.A1(_00438_),
    .A2(_01724_),
    .A3(_01649_),
    .ZN(_01725_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _07336_ (.A1(_01564_),
    .A2(_01565_),
    .A3(_01648_),
    .B(_01725_),
    .ZN(_01726_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07337_ (.A1(_01658_),
    .A2(_01662_),
    .ZN(_01727_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07338_ (.A1(_01653_),
    .A2(_01727_),
    .ZN(_01728_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _07339_ (.A1(_01651_),
    .A2(_01663_),
    .B(_01728_),
    .ZN(_01729_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07340_ (.A1(_01656_),
    .A2(_01657_),
    .ZN(_01730_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07341_ (.A1(_01656_),
    .A2(_01657_),
    .ZN(_01731_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07342_ (.A1(_01655_),
    .A2(_01730_),
    .B(_01731_),
    .ZN(_01732_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07343_ (.I(_01557_),
    .Z(_01733_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07344_ (.A1(_05817_),
    .A2(_01733_),
    .ZN(_01734_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07345_ (.A1(_01732_),
    .A2(_01734_),
    .ZN(_01735_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07346_ (.A1(_05808_),
    .A2(_01467_),
    .ZN(_01736_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07347_ (.A1(_01735_),
    .A2(_01736_),
    .Z(_01737_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _07348_ (.A1(_05796_),
    .A2(_05806_),
    .A3(_01390_),
    .A4(_01386_),
    .Z(_01738_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07349_ (.A1(_01568_),
    .A2(_01738_),
    .ZN(_01739_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07350_ (.A1(_01658_),
    .A2(_01659_),
    .A3(_01661_),
    .ZN(_01740_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07351_ (.A1(_01739_),
    .A2(_01740_),
    .ZN(_01741_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07352_ (.I(_01654_),
    .Z(_01742_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07353_ (.A1(_01383_),
    .A2(_01742_),
    .Z(_01743_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07354_ (.A1(_05854_),
    .A2(_01472_),
    .ZN(_01744_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07355_ (.A1(_05757_),
    .A2(_01144_),
    .ZN(_01745_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _07356_ (.A1(_01743_),
    .A2(_01744_),
    .A3(_01745_),
    .ZN(_01746_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07357_ (.A1(\as2650.r0[5] ),
    .A2(_01310_),
    .ZN(_01747_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07358_ (.A1(\as2650.r0[4] ),
    .A2(_01384_),
    .ZN(_01748_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07359_ (.A1(\as2650.r0[0] ),
    .A2(_05765_),
    .ZN(_01749_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _07360_ (.A1(_01747_),
    .A2(_01748_),
    .A3(_01749_),
    .Z(_01750_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07361_ (.A1(_01738_),
    .A2(_01750_),
    .Z(_01751_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07362_ (.A1(_01746_),
    .A2(_01751_),
    .ZN(_01752_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07363_ (.A1(_01741_),
    .A2(_01752_),
    .Z(_01753_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07364_ (.A1(_01737_),
    .A2(_01753_),
    .Z(_01754_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07365_ (.A1(_01729_),
    .A2(_01754_),
    .Z(_01755_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07366_ (.A1(_01726_),
    .A2(_01755_),
    .Z(_01756_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07367_ (.A1(_01723_),
    .A2(_01756_),
    .ZN(_01757_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _07368_ (.A1(_01720_),
    .A2(_01757_),
    .ZN(_01758_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07369_ (.A1(\as2650.r123[1][7] ),
    .A2(_01154_),
    .ZN(_01759_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _07370_ (.A1(_01046_),
    .A2(_01718_),
    .B1(_01758_),
    .B2(_01403_),
    .C(_01759_),
    .ZN(_00021_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07371_ (.I(_01132_),
    .Z(_01760_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07372_ (.I(_01760_),
    .Z(_01761_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07373_ (.I(_01761_),
    .Z(_01762_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07374_ (.I(_01001_),
    .Z(_01763_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _07375_ (.A1(_00821_),
    .A2(_00955_),
    .ZN(_01764_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07376_ (.A1(_00836_),
    .A2(_01763_),
    .A3(_01764_),
    .ZN(_01765_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07377_ (.I(_01765_),
    .Z(_01766_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07378_ (.I(_01766_),
    .Z(_01767_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07379_ (.I(net59),
    .ZN(_01768_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07380_ (.I(_01768_),
    .Z(_01769_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _07381_ (.I(net90),
    .ZN(_01770_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _07382_ (.A1(_01769_),
    .A2(_01770_),
    .ZN(_01771_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07383_ (.I(_01771_),
    .Z(_01772_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07384_ (.I(net70),
    .Z(_01773_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07385_ (.I(_01773_),
    .Z(_01774_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07386_ (.I(_01774_),
    .Z(_01775_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07387_ (.I(net73),
    .Z(_01776_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07388_ (.I(_01776_),
    .Z(_01777_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07389_ (.A1(_01775_),
    .A2(_01777_),
    .ZN(_01778_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07390_ (.I(_01778_),
    .Z(_01779_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07391_ (.A1(_01767_),
    .A2(_01772_),
    .A3(_01779_),
    .ZN(_01780_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07392_ (.I(_01780_),
    .Z(_01781_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07393_ (.I(_01781_),
    .Z(_01782_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07394_ (.I(_01775_),
    .Z(_01783_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07395_ (.I(_01777_),
    .Z(_01784_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07396_ (.I(_01784_),
    .Z(_01785_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07397_ (.I(_01765_),
    .ZN(_01786_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _07398_ (.A1(_00971_),
    .A2(_00973_),
    .Z(_01787_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _07399_ (.A1(_01787_),
    .A2(_01022_),
    .Z(_01788_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07400_ (.A1(_01786_),
    .A2(_01788_),
    .ZN(_01789_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _07401_ (.A1(_00689_),
    .A2(\as2650.last_intr ),
    .A3(net75),
    .Z(_01790_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _07402_ (.A1(_00515_),
    .A2(_01790_),
    .ZN(_01791_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _07403_ (.A1(_00578_),
    .A2(_01791_),
    .ZN(_01792_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07404_ (.A1(\as2650.cycle[6] ),
    .A2(_00643_),
    .ZN(_01793_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07405_ (.A1(_00509_),
    .A2(net3),
    .ZN(_01794_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07406_ (.A1(_00757_),
    .A2(_00915_),
    .ZN(_01795_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07407_ (.A1(_00889_),
    .A2(_01795_),
    .B(_00579_),
    .ZN(_01796_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07408_ (.A1(_01793_),
    .A2(_01794_),
    .B1(_01796_),
    .B2(_00864_),
    .ZN(_01797_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07409_ (.A1(_00549_),
    .A2(_00874_),
    .ZN(_01798_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _07410_ (.A1(_05740_),
    .A2(_05756_),
    .B(_00500_),
    .ZN(_01799_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07411_ (.A1(_01798_),
    .A2(_01799_),
    .ZN(_01800_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07412_ (.A1(_00683_),
    .A2(_00737_),
    .ZN(_01801_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07413_ (.I(_01016_),
    .Z(_01802_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07414_ (.A1(_01802_),
    .A2(_00697_),
    .A3(_00674_),
    .ZN(_01803_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _07415_ (.A1(_00540_),
    .A2(_01797_),
    .A3(_01800_),
    .B1(_01801_),
    .B2(_01803_),
    .ZN(_01804_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07416_ (.A1(_01763_),
    .A2(_01804_),
    .ZN(_01805_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07417_ (.A1(_01789_),
    .A2(_01792_),
    .A3(_01805_),
    .ZN(_01806_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07418_ (.I(_01806_),
    .Z(_01807_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07419_ (.I(net59),
    .Z(_01808_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07420_ (.A1(_01808_),
    .A2(_01770_),
    .ZN(_01809_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07421_ (.I(_01809_),
    .Z(_01810_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07422_ (.I(_01810_),
    .Z(_01811_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07423_ (.I(_01811_),
    .Z(_01812_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07424_ (.I(_01812_),
    .Z(_01813_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07425_ (.I(_01813_),
    .Z(_01814_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07426_ (.I(_01814_),
    .Z(_01815_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07427_ (.I(_01815_),
    .Z(_01816_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _07428_ (.A1(_01783_),
    .A2(_01785_),
    .A3(_01807_),
    .A4(_01816_),
    .ZN(_01817_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07429_ (.I(_01817_),
    .Z(_01818_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07430_ (.A1(\as2650.stack[13][0] ),
    .A2(_01818_),
    .ZN(_01819_));
 gf180mcu_fd_sc_mcu7t5v0__and3_2 _07431_ (.A1(_01789_),
    .A2(_01792_),
    .A3(_01805_),
    .Z(_01820_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07432_ (.I(_01820_),
    .Z(_01821_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07433_ (.I(_01769_),
    .Z(_01822_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07434_ (.I(net90),
    .Z(_01823_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07435_ (.A1(_01822_),
    .A2(_01823_),
    .ZN(_01824_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _07436_ (.I(_01824_),
    .Z(_01825_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _07437_ (.A1(_01779_),
    .A2(_01821_),
    .A3(_01825_),
    .ZN(_01826_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07438_ (.I(_01826_),
    .Z(_01827_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07439_ (.I(_01827_),
    .Z(_01828_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07440_ (.I(_01053_),
    .ZN(_01829_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07441_ (.I(_01829_),
    .Z(_01830_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07442_ (.I(_01789_),
    .Z(_01831_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07443_ (.I(_01831_),
    .Z(_01832_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07444_ (.I(_01832_),
    .Z(_01833_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07445_ (.I(net55),
    .Z(_01834_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07446_ (.I(_01834_),
    .Z(_01835_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07447_ (.I(_01835_),
    .Z(_01836_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07448_ (.I(_01831_),
    .Z(_01837_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _07449_ (.A1(_01836_),
    .A2(_01837_),
    .ZN(_01838_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _07450_ (.A1(_01830_),
    .A2(_01833_),
    .B(_01838_),
    .ZN(_01839_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07451_ (.I(_01839_),
    .Z(_01840_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07452_ (.I(_01780_),
    .Z(_01841_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07453_ (.I(_01841_),
    .Z(_01842_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _07454_ (.A1(_01828_),
    .A2(_01840_),
    .B(_01842_),
    .ZN(_01843_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07455_ (.A1(_01762_),
    .A2(_01782_),
    .B1(_01819_),
    .B2(_01843_),
    .ZN(_00022_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07456_ (.I(net79),
    .ZN(_01844_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07457_ (.I(_01844_),
    .Z(_01845_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07458_ (.I(_01845_),
    .Z(_01846_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07459_ (.I(_01846_),
    .Z(_01847_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07460_ (.A1(\as2650.stack[13][1] ),
    .A2(_01818_),
    .ZN(_01848_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07461_ (.I(_01826_),
    .Z(_01849_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07462_ (.I(_01209_),
    .Z(_01850_));
 gf180mcu_fd_sc_mcu7t5v0__inv_4 _07463_ (.I(_01850_),
    .ZN(_01851_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07464_ (.I(_01831_),
    .Z(_01852_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07465_ (.I(net56),
    .Z(_01853_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07466_ (.I(_01853_),
    .Z(_01854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07467_ (.I(_01854_),
    .Z(_01855_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07468_ (.A1(_01855_),
    .A2(_01837_),
    .ZN(_01856_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _07469_ (.A1(_01851_),
    .A2(_01852_),
    .B(_01856_),
    .ZN(_01857_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07470_ (.I(_01857_),
    .Z(_01858_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07471_ (.I(_01841_),
    .Z(_01859_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07472_ (.A1(_01849_),
    .A2(_01858_),
    .B(_01859_),
    .ZN(_01860_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07473_ (.A1(_01847_),
    .A2(_01782_),
    .B1(_01848_),
    .B2(_01860_),
    .ZN(_00023_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _07474_ (.I(net49),
    .ZN(_01861_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07475_ (.I(_01861_),
    .Z(_01862_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07476_ (.I(_01862_),
    .Z(_01863_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07477_ (.A1(\as2650.stack[13][2] ),
    .A2(_01818_),
    .ZN(_01864_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07478_ (.I(_01272_),
    .Z(_01865_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07479_ (.I(net57),
    .Z(_01866_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07480_ (.I(_01866_),
    .Z(_01867_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07481_ (.I(_01867_),
    .Z(_01868_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07482_ (.I0(_01865_),
    .I1(_01868_),
    .S(_01832_),
    .Z(_01869_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07483_ (.I(_01869_),
    .Z(_01870_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07484_ (.A1(_01849_),
    .A2(_01870_),
    .B(_01859_),
    .ZN(_01871_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07485_ (.A1(_01863_),
    .A2(_01782_),
    .B1(_01864_),
    .B2(_01871_),
    .ZN(_00024_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _07486_ (.I(_01065_),
    .ZN(_01872_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07487_ (.I(_01872_),
    .Z(_01873_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07488_ (.I(_01873_),
    .Z(_01874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07489_ (.A1(\as2650.stack[13][3] ),
    .A2(_01818_),
    .ZN(_01875_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07490_ (.I(net58),
    .ZN(_01876_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07491_ (.I(_01876_),
    .Z(_01877_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07492_ (.I(_01831_),
    .Z(_01878_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07493_ (.A1(_01325_),
    .A2(_01878_),
    .ZN(_01879_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _07494_ (.A1(_01877_),
    .A2(_01837_),
    .B(_01879_),
    .ZN(_01880_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07495_ (.I(_01880_),
    .Z(_01881_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07496_ (.A1(_01849_),
    .A2(_01881_),
    .B(_01859_),
    .ZN(_01882_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07497_ (.A1(_01874_),
    .A2(_01782_),
    .B1(_01875_),
    .B2(_01882_),
    .ZN(_00025_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07498_ (.I(_01147_),
    .Z(_01883_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07499_ (.I(_01883_),
    .Z(_01884_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07500_ (.I(_01841_),
    .Z(_01885_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07501_ (.I(_01817_),
    .Z(_01886_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07502_ (.A1(\as2650.stack[13][4] ),
    .A2(_01886_),
    .ZN(_01887_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07503_ (.I(net60),
    .ZN(_01888_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07504_ (.I(_01888_),
    .Z(_01889_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07505_ (.A1(_01421_),
    .A2(_01832_),
    .ZN(_01890_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _07506_ (.A1(_01889_),
    .A2(_01837_),
    .B(_01890_),
    .ZN(_01891_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07507_ (.I(_01891_),
    .Z(_01892_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07508_ (.A1(_01849_),
    .A2(_01892_),
    .B(_01859_),
    .ZN(_01893_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07509_ (.A1(_01884_),
    .A2(_01885_),
    .B1(_01887_),
    .B2(_01893_),
    .ZN(_00026_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07510_ (.I(net52),
    .ZN(_01894_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07511_ (.I(_01894_),
    .Z(_01895_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07512_ (.I(_01895_),
    .Z(_01896_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07513_ (.A1(\as2650.stack[13][5] ),
    .A2(_01886_),
    .ZN(_01897_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07514_ (.I(_01826_),
    .Z(_01898_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _07515_ (.I(_01533_),
    .ZN(_01899_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07516_ (.I(_01899_),
    .Z(_01900_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07517_ (.I(net61),
    .Z(_01901_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07518_ (.I(_01901_),
    .Z(_01902_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07519_ (.I(_01902_),
    .Z(_01903_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07520_ (.A1(_01903_),
    .A2(_01878_),
    .ZN(_01904_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _07521_ (.A1(_01900_),
    .A2(_01852_),
    .B(_01904_),
    .ZN(_01905_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07522_ (.I(_01905_),
    .Z(_01906_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07523_ (.A1(_01898_),
    .A2(_01906_),
    .B(_01781_),
    .ZN(_01907_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07524_ (.A1(_01896_),
    .A2(_01885_),
    .B1(_01897_),
    .B2(_01907_),
    .ZN(_00027_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07525_ (.I(_05735_),
    .Z(_01908_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07526_ (.I(_01908_),
    .Z(_01909_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07527_ (.A1(\as2650.stack[13][6] ),
    .A2(_01886_),
    .ZN(_01910_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _07528_ (.I(_01615_),
    .ZN(_01911_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07529_ (.I(net62),
    .Z(_01912_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07530_ (.I(_01912_),
    .Z(_01913_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07531_ (.A1(_01913_),
    .A2(_01878_),
    .ZN(_01914_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07532_ (.A1(_01911_),
    .A2(_01852_),
    .B(_01914_),
    .ZN(_01915_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07533_ (.I(_01915_),
    .Z(_01916_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07534_ (.A1(_01898_),
    .A2(_01916_),
    .B(_01781_),
    .ZN(_01917_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07535_ (.A1(_01909_),
    .A2(_01885_),
    .B1(_01910_),
    .B2(_01917_),
    .ZN(_00028_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07536_ (.I(_05727_),
    .Z(_01918_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07537_ (.I(_01918_),
    .Z(_01919_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07538_ (.A1(\as2650.stack[13][7] ),
    .A2(_01886_),
    .ZN(_01920_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _07539_ (.I(_01674_),
    .ZN(_01921_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07540_ (.I(net93),
    .Z(_01922_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _07541_ (.A1(_01922_),
    .A2(_01878_),
    .ZN(_01923_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _07542_ (.A1(_01921_),
    .A2(_01852_),
    .B(_01923_),
    .ZN(_01924_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07543_ (.I(_01924_),
    .Z(_01925_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07544_ (.A1(_01898_),
    .A2(_01925_),
    .B(_01781_),
    .ZN(_01926_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07545_ (.A1(_01919_),
    .A2(_01885_),
    .B1(_01920_),
    .B2(_01926_),
    .ZN(_00029_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07546_ (.A1(_00901_),
    .A2(_00980_),
    .A3(_00964_),
    .ZN(_01927_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07547_ (.I(_01927_),
    .Z(_01928_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07548_ (.I(_01928_),
    .Z(_01929_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07549_ (.I(_01929_),
    .Z(_01930_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07550_ (.A1(_01930_),
    .A2(_00984_),
    .B(_01149_),
    .ZN(_01931_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07551_ (.A1(_01150_),
    .A2(_01931_),
    .ZN(_01932_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07552_ (.I(_01932_),
    .Z(_01933_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _07553_ (.A1(_01147_),
    .A2(_00942_),
    .A3(_01400_),
    .ZN(_01934_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07554_ (.I(_01934_),
    .Z(_01935_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _07555_ (.I(net70),
    .ZN(_01936_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07556_ (.A1(_01936_),
    .A2(net73),
    .ZN(_01937_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07557_ (.A1(_01771_),
    .A2(_01937_),
    .ZN(_01938_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07558_ (.A1(net59),
    .A2(net90),
    .ZN(_01939_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07559_ (.I(_01939_),
    .Z(_01940_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07560_ (.A1(_01936_),
    .A2(_01940_),
    .B(net73),
    .ZN(_01941_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07561_ (.A1(_01938_),
    .A2(_01941_),
    .ZN(_01942_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07562_ (.I(_01942_),
    .Z(_01943_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07563_ (.I(_01943_),
    .Z(_01944_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07564_ (.I(_01944_),
    .Z(_01945_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _07565_ (.A1(net70),
    .A2(_01939_),
    .Z(_01946_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _07566_ (.I(_01946_),
    .ZN(_01947_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07567_ (.I(_01947_),
    .Z(_01948_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07568_ (.I(_01948_),
    .Z(_01949_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07569_ (.I(_01949_),
    .Z(_01950_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07570_ (.I(_01812_),
    .Z(_01951_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07571_ (.A1(_01768_),
    .A2(net48),
    .ZN(_01952_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07572_ (.I(_01952_),
    .Z(_01953_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07573_ (.I(_01953_),
    .Z(_01954_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07574_ (.I(_01954_),
    .Z(_01955_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07575_ (.I(_01955_),
    .Z(_01956_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07576_ (.A1(\as2650.stack[8][8] ),
    .A2(_01951_),
    .B1(_01956_),
    .B2(\as2650.stack[9][8] ),
    .ZN(_01957_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07577_ (.I(_01939_),
    .Z(_01958_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07578_ (.I(_01958_),
    .Z(_01959_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07579_ (.I(_01959_),
    .Z(_01960_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07580_ (.I(_01960_),
    .Z(_01961_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07581_ (.A1(_01768_),
    .A2(_01770_),
    .ZN(_01962_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07582_ (.I(_01962_),
    .Z(_01963_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07583_ (.I(_01963_),
    .Z(_01964_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07584_ (.I(_01964_),
    .Z(_01965_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07585_ (.I(_01965_),
    .Z(_01966_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07586_ (.A1(\as2650.stack[11][8] ),
    .A2(_01961_),
    .B1(_01966_),
    .B2(\as2650.stack[10][8] ),
    .ZN(_01967_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07587_ (.A1(_01950_),
    .A2(_01957_),
    .A3(_01967_),
    .ZN(_01968_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07588_ (.I(_01946_),
    .Z(_01969_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07589_ (.I(_01969_),
    .Z(_01970_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07590_ (.I(_01970_),
    .Z(_01971_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07591_ (.A1(\as2650.stack[15][8] ),
    .A2(_01961_),
    .B1(_01966_),
    .B2(\as2650.stack[14][8] ),
    .ZN(_01972_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07592_ (.A1(\as2650.stack[12][8] ),
    .A2(_01951_),
    .B1(_01956_),
    .B2(\as2650.stack[13][8] ),
    .ZN(_01973_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07593_ (.A1(_01971_),
    .A2(_01972_),
    .A3(_01973_),
    .ZN(_01974_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07594_ (.A1(_01968_),
    .A2(_01974_),
    .ZN(_01975_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07595_ (.I(_01812_),
    .Z(_01976_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07596_ (.I(_01955_),
    .Z(_01977_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07597_ (.A1(\as2650.stack[0][8] ),
    .A2(_01976_),
    .B1(_01977_),
    .B2(\as2650.stack[1][8] ),
    .ZN(_01978_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07598_ (.I(_01940_),
    .Z(_01979_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07599_ (.I(_01979_),
    .Z(_01980_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07600_ (.I(_01980_),
    .Z(_01981_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07601_ (.I(_01965_),
    .Z(_01982_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07602_ (.A1(\as2650.stack[3][8] ),
    .A2(_01981_),
    .B1(_01982_),
    .B2(\as2650.stack[2][8] ),
    .ZN(_01983_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07603_ (.A1(_01950_),
    .A2(_01978_),
    .A3(_01983_),
    .ZN(_01984_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07604_ (.I(_01980_),
    .Z(_01985_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07605_ (.A1(\as2650.stack[7][8] ),
    .A2(_01985_),
    .B1(_01982_),
    .B2(\as2650.stack[6][8] ),
    .ZN(_01986_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07606_ (.A1(\as2650.stack[4][8] ),
    .A2(_01976_),
    .B1(_01977_),
    .B2(\as2650.stack[5][8] ),
    .ZN(_01987_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07607_ (.A1(_01971_),
    .A2(_01986_),
    .A3(_01987_),
    .ZN(_01988_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07608_ (.A1(_01984_),
    .A2(_01988_),
    .B(_01945_),
    .ZN(_01989_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _07609_ (.A1(_01945_),
    .A2(_01975_),
    .B(_01989_),
    .ZN(_01990_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07610_ (.A1(_01935_),
    .A2(_01990_),
    .ZN(_01991_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07611_ (.A1(_01930_),
    .A2(_01149_),
    .ZN(_01992_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07612_ (.I(_01992_),
    .Z(_01993_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07613_ (.A1(_01142_),
    .A2(_01993_),
    .ZN(_01994_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07614_ (.A1(_05763_),
    .A2(_01043_),
    .ZN(_01995_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07615_ (.I(_01995_),
    .Z(_01996_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _07616_ (.A1(_01933_),
    .A2(_01991_),
    .A3(_01994_),
    .B1(_01996_),
    .B2(_01141_),
    .ZN(_01997_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07617_ (.A1(_05718_),
    .A2(_01931_),
    .ZN(_01998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07618_ (.A1(_01995_),
    .A2(_01998_),
    .ZN(_01999_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07619_ (.I(_01999_),
    .Z(_02000_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07620_ (.I0(\as2650.r123[0][0] ),
    .I1(_01997_),
    .S(_02000_),
    .Z(_02001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07621_ (.I(_02001_),
    .Z(_00030_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07622_ (.I(_01945_),
    .Z(_02002_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07623_ (.I(_01950_),
    .Z(_02003_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07624_ (.I(_01951_),
    .Z(_02004_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07625_ (.I(_01956_),
    .Z(_02005_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07626_ (.A1(\as2650.stack[8][9] ),
    .A2(_02004_),
    .B1(_02005_),
    .B2(\as2650.stack[9][9] ),
    .ZN(_02006_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07627_ (.I(_01981_),
    .Z(_02007_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07628_ (.I(_01966_),
    .Z(_02008_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07629_ (.A1(\as2650.stack[11][9] ),
    .A2(_02007_),
    .B1(_02008_),
    .B2(\as2650.stack[10][9] ),
    .ZN(_02009_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07630_ (.A1(_02003_),
    .A2(_02006_),
    .A3(_02009_),
    .ZN(_02010_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07631_ (.I(_01971_),
    .Z(_02011_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07632_ (.I(_01981_),
    .Z(_02012_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07633_ (.I(_01982_),
    .Z(_02013_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07634_ (.A1(\as2650.stack[15][9] ),
    .A2(_02012_),
    .B1(_02013_),
    .B2(\as2650.stack[14][9] ),
    .ZN(_02014_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07635_ (.I(_01976_),
    .Z(_02015_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07636_ (.I(_01977_),
    .Z(_02016_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07637_ (.A1(\as2650.stack[12][9] ),
    .A2(_02015_),
    .B1(_02016_),
    .B2(\as2650.stack[13][9] ),
    .ZN(_02017_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07638_ (.A1(_02011_),
    .A2(_02014_),
    .A3(_02017_),
    .ZN(_02018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07639_ (.A1(_02010_),
    .A2(_02018_),
    .ZN(_02019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07640_ (.I(_01949_),
    .Z(_02020_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07641_ (.I(_01976_),
    .Z(_02021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07642_ (.I(_01977_),
    .Z(_02022_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07643_ (.A1(\as2650.stack[0][9] ),
    .A2(_02021_),
    .B1(_02022_),
    .B2(\as2650.stack[1][9] ),
    .ZN(_02023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07644_ (.I(_01985_),
    .Z(_02024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07645_ (.I(_01982_),
    .Z(_02025_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07646_ (.A1(\as2650.stack[3][9] ),
    .A2(_02024_),
    .B1(_02025_),
    .B2(\as2650.stack[2][9] ),
    .ZN(_02026_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07647_ (.A1(_02020_),
    .A2(_02023_),
    .A3(_02026_),
    .ZN(_02027_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07648_ (.I(_01971_),
    .Z(_02028_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07649_ (.I(_01985_),
    .Z(_02029_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07650_ (.I(_01962_),
    .Z(_02030_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07651_ (.I(_02030_),
    .Z(_02031_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07652_ (.I(_02031_),
    .Z(_02032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07653_ (.I(_02032_),
    .Z(_02033_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07654_ (.A1(\as2650.stack[7][9] ),
    .A2(_02029_),
    .B1(_02033_),
    .B2(\as2650.stack[6][9] ),
    .ZN(_02034_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07655_ (.I(_01813_),
    .Z(_02035_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07656_ (.I(_01955_),
    .Z(_02036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07657_ (.I(_02036_),
    .Z(_02037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _07658_ (.A1(\as2650.stack[4][9] ),
    .A2(_02035_),
    .B1(_02037_),
    .B2(\as2650.stack[5][9] ),
    .ZN(_02038_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07659_ (.A1(_02028_),
    .A2(_02034_),
    .A3(_02038_),
    .ZN(_02039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07660_ (.I(_01944_),
    .Z(_02040_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07661_ (.A1(_02027_),
    .A2(_02039_),
    .B(_02040_),
    .ZN(_02041_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _07662_ (.A1(_02002_),
    .A2(_02019_),
    .B(_02041_),
    .ZN(_02042_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07663_ (.A1(_01935_),
    .A2(_02042_),
    .ZN(_02043_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07664_ (.A1(_01850_),
    .A2(_01993_),
    .ZN(_02044_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _07665_ (.A1(_01933_),
    .A2(_02043_),
    .A3(_02044_),
    .B1(_01996_),
    .B2(_01233_),
    .ZN(_02045_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07666_ (.I0(\as2650.r123[0][1] ),
    .I1(_02045_),
    .S(_02000_),
    .Z(_02046_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07667_ (.I(_02046_),
    .Z(_00031_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07668_ (.A1(\as2650.stack[8][10] ),
    .A2(_02004_),
    .B1(_02005_),
    .B2(\as2650.stack[9][10] ),
    .ZN(_02047_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07669_ (.A1(\as2650.stack[11][10] ),
    .A2(_02007_),
    .B1(_02008_),
    .B2(\as2650.stack[10][10] ),
    .ZN(_02048_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07670_ (.A1(_02003_),
    .A2(_02047_),
    .A3(_02048_),
    .ZN(_02049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07671_ (.A1(\as2650.stack[15][10] ),
    .A2(_02012_),
    .B1(_02013_),
    .B2(\as2650.stack[14][10] ),
    .ZN(_02050_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07672_ (.A1(\as2650.stack[12][10] ),
    .A2(_02015_),
    .B1(_02016_),
    .B2(\as2650.stack[13][10] ),
    .ZN(_02051_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07673_ (.A1(_02011_),
    .A2(_02050_),
    .A3(_02051_),
    .ZN(_02052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07674_ (.A1(_02049_),
    .A2(_02052_),
    .ZN(_02053_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07675_ (.I(_01813_),
    .Z(_02054_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07676_ (.A1(\as2650.stack[0][10] ),
    .A2(_02054_),
    .B1(_02022_),
    .B2(\as2650.stack[1][10] ),
    .ZN(_02055_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07677_ (.I(_02032_),
    .Z(_02056_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07678_ (.A1(\as2650.stack[3][10] ),
    .A2(_02024_),
    .B1(_02056_),
    .B2(\as2650.stack[2][10] ),
    .ZN(_02057_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07679_ (.A1(_02020_),
    .A2(_02055_),
    .A3(_02057_),
    .ZN(_02058_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07680_ (.I(_01985_),
    .Z(_02059_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07681_ (.A1(\as2650.stack[7][10] ),
    .A2(_02059_),
    .B1(_02033_),
    .B2(\as2650.stack[6][10] ),
    .ZN(_02060_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07682_ (.I(_02036_),
    .Z(_02061_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _07683_ (.A1(\as2650.stack[4][10] ),
    .A2(_02035_),
    .B1(_02061_),
    .B2(\as2650.stack[5][10] ),
    .ZN(_02062_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07684_ (.A1(_02028_),
    .A2(_02060_),
    .A3(_02062_),
    .ZN(_02063_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07685_ (.A1(_02058_),
    .A2(_02063_),
    .B(_02040_),
    .ZN(_02064_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _07686_ (.A1(_02002_),
    .A2(_02053_),
    .B(_02064_),
    .ZN(_02065_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07687_ (.A1(_01935_),
    .A2(_02065_),
    .ZN(_02066_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07688_ (.I(_01272_),
    .Z(_02067_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07689_ (.A1(_02067_),
    .A2(_01993_),
    .ZN(_02068_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _07690_ (.A1(_01933_),
    .A2(_02066_),
    .A3(_02068_),
    .B1(_01996_),
    .B2(_01305_),
    .ZN(_02069_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07691_ (.I0(\as2650.r123[0][2] ),
    .I1(_02069_),
    .S(_02000_),
    .Z(_02070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07692_ (.I(_02070_),
    .Z(_00032_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07693_ (.I(_01932_),
    .Z(_02071_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07694_ (.A1(\as2650.stack[8][11] ),
    .A2(_02021_),
    .B1(_02022_),
    .B2(\as2650.stack[9][11] ),
    .ZN(_02072_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07695_ (.A1(\as2650.stack[11][11] ),
    .A2(_02024_),
    .B1(_02025_),
    .B2(\as2650.stack[10][11] ),
    .ZN(_02073_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07696_ (.A1(_02020_),
    .A2(_02072_),
    .A3(_02073_),
    .ZN(_02074_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07697_ (.A1(\as2650.stack[15][11] ),
    .A2(_02024_),
    .B1(_02025_),
    .B2(\as2650.stack[14][11] ),
    .ZN(_02075_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07698_ (.A1(\as2650.stack[12][11] ),
    .A2(_02021_),
    .B1(_02022_),
    .B2(\as2650.stack[13][11] ),
    .ZN(_02076_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07699_ (.A1(_02011_),
    .A2(_02075_),
    .A3(_02076_),
    .ZN(_02077_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07700_ (.A1(_02074_),
    .A2(_02077_),
    .ZN(_02078_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07701_ (.I(_01949_),
    .Z(_02079_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07702_ (.I(_02036_),
    .Z(_02080_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07703_ (.A1(\as2650.stack[0][11] ),
    .A2(_01814_),
    .B1(_02080_),
    .B2(\as2650.stack[1][11] ),
    .ZN(_02081_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07704_ (.I(_01960_),
    .Z(_02082_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07705_ (.I(_02032_),
    .Z(_02083_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07706_ (.A1(\as2650.stack[3][11] ),
    .A2(_02082_),
    .B1(_02083_),
    .B2(\as2650.stack[2][11] ),
    .ZN(_02084_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07707_ (.A1(_02079_),
    .A2(_02081_),
    .A3(_02084_),
    .ZN(_02085_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07708_ (.I(_01970_),
    .Z(_02086_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07709_ (.I(_01960_),
    .Z(_02087_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07710_ (.A1(\as2650.stack[7][11] ),
    .A2(_02087_),
    .B1(_02083_),
    .B2(\as2650.stack[6][11] ),
    .ZN(_02088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07711_ (.I(_01813_),
    .Z(_02089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07712_ (.I(_02036_),
    .Z(_02090_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07713_ (.A1(\as2650.stack[4][11] ),
    .A2(_02089_),
    .B1(_02090_),
    .B2(\as2650.stack[5][11] ),
    .ZN(_02091_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07714_ (.A1(_02086_),
    .A2(_02088_),
    .A3(_02091_),
    .ZN(_02092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07715_ (.I(_01944_),
    .Z(_02093_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07716_ (.A1(_02085_),
    .A2(_02092_),
    .B(_02093_),
    .ZN(_02094_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _07717_ (.A1(_02002_),
    .A2(_02078_),
    .B(_02094_),
    .ZN(_02095_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07718_ (.A1(_01935_),
    .A2(_02095_),
    .ZN(_02096_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07719_ (.I(_01325_),
    .Z(_02097_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07720_ (.I(_02097_),
    .Z(_02098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07721_ (.I(_01992_),
    .Z(_02099_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07722_ (.A1(_02098_),
    .A2(_02099_),
    .ZN(_02100_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07723_ (.I(_01995_),
    .Z(_02101_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _07724_ (.A1(_02071_),
    .A2(_02096_),
    .A3(_02100_),
    .B1(_02101_),
    .B2(_01375_),
    .ZN(_02102_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07725_ (.I0(\as2650.r123[0][3] ),
    .I1(_02102_),
    .S(_02000_),
    .Z(_02103_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07726_ (.I(_02103_),
    .Z(_00033_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07727_ (.A1(\as2650.stack[8][12] ),
    .A2(_02015_),
    .B1(_02005_),
    .B2(\as2650.stack[9][12] ),
    .ZN(_02104_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07728_ (.A1(\as2650.stack[11][12] ),
    .A2(_02012_),
    .B1(_02008_),
    .B2(\as2650.stack[10][12] ),
    .ZN(_02105_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07729_ (.A1(_02003_),
    .A2(_02104_),
    .A3(_02105_),
    .ZN(_02106_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07730_ (.A1(\as2650.stack[15][12] ),
    .A2(_02012_),
    .B1(_02013_),
    .B2(\as2650.stack[14][12] ),
    .ZN(_02107_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07731_ (.A1(\as2650.stack[12][12] ),
    .A2(_02015_),
    .B1(_02016_),
    .B2(\as2650.stack[13][12] ),
    .ZN(_02108_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07732_ (.A1(_02011_),
    .A2(_02107_),
    .A3(_02108_),
    .ZN(_02109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _07733_ (.A1(_02106_),
    .A2(_02109_),
    .ZN(_02110_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07734_ (.A1(\as2650.stack[0][12] ),
    .A2(_02054_),
    .B1(_02037_),
    .B2(\as2650.stack[1][12] ),
    .ZN(_02111_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07735_ (.A1(\as2650.stack[3][12] ),
    .A2(_02029_),
    .B1(_02056_),
    .B2(\as2650.stack[2][12] ),
    .ZN(_02112_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07736_ (.A1(_02020_),
    .A2(_02111_),
    .A3(_02112_),
    .ZN(_02113_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07737_ (.A1(\as2650.stack[7][12] ),
    .A2(_02059_),
    .B1(_02033_),
    .B2(\as2650.stack[6][12] ),
    .ZN(_02114_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07738_ (.A1(\as2650.stack[4][12] ),
    .A2(_02035_),
    .B1(_02061_),
    .B2(\as2650.stack[5][12] ),
    .ZN(_02115_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07739_ (.A1(_02028_),
    .A2(_02114_),
    .A3(_02115_),
    .ZN(_02116_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07740_ (.A1(_02113_),
    .A2(_02116_),
    .B(_02093_),
    .ZN(_02117_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _07741_ (.A1(_02002_),
    .A2(_02110_),
    .B(_02117_),
    .ZN(_02118_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07742_ (.A1(_01934_),
    .A2(_02118_),
    .ZN(_02119_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07743_ (.I(_01421_),
    .Z(_02120_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07744_ (.A1(_02120_),
    .A2(_02099_),
    .ZN(_02121_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _07745_ (.A1(_02071_),
    .A2(_02119_),
    .A3(_02121_),
    .B1(_02101_),
    .B2(_01462_),
    .ZN(_02122_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07746_ (.I(_01999_),
    .Z(_02123_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07747_ (.I0(\as2650.r123[0][4] ),
    .I1(_02122_),
    .S(_02123_),
    .Z(_02124_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07748_ (.I(_02124_),
    .Z(_00034_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07749_ (.A1(\as2650.stack[8][13] ),
    .A2(_02089_),
    .B1(_02090_),
    .B2(\as2650.stack[9][13] ),
    .ZN(_02125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07750_ (.I(_02032_),
    .Z(_02126_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07751_ (.A1(\as2650.stack[11][13] ),
    .A2(_02087_),
    .B1(_02126_),
    .B2(\as2650.stack[10][13] ),
    .ZN(_02127_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07752_ (.A1(_02079_),
    .A2(_02125_),
    .A3(_02127_),
    .ZN(_02128_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07753_ (.I(_01960_),
    .Z(_02129_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07754_ (.A1(\as2650.stack[15][13] ),
    .A2(_02129_),
    .B1(_02126_),
    .B2(\as2650.stack[14][13] ),
    .ZN(_02130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07755_ (.I(_01812_),
    .Z(_02131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07756_ (.I(_01955_),
    .Z(_02132_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07757_ (.A1(\as2650.stack[12][13] ),
    .A2(_02131_),
    .B1(_02132_),
    .B2(\as2650.stack[13][13] ),
    .ZN(_02133_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07758_ (.A1(_02086_),
    .A2(_02130_),
    .A3(_02133_),
    .ZN(_02134_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07759_ (.A1(_02128_),
    .A2(_02134_),
    .ZN(_02135_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07760_ (.A1(\as2650.stack[0][13] ),
    .A2(_02131_),
    .B1(_02132_),
    .B2(\as2650.stack[1][13] ),
    .ZN(_02136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07761_ (.I(_01965_),
    .Z(_02137_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07762_ (.A1(\as2650.stack[3][13] ),
    .A2(_02129_),
    .B1(_02137_),
    .B2(\as2650.stack[2][13] ),
    .ZN(_02138_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07763_ (.A1(_01950_),
    .A2(_02136_),
    .A3(_02138_),
    .ZN(_02139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07764_ (.A1(\as2650.stack[7][13] ),
    .A2(_01961_),
    .B1(_02137_),
    .B2(\as2650.stack[6][13] ),
    .ZN(_02140_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07765_ (.A1(\as2650.stack[4][13] ),
    .A2(_01951_),
    .B1(_01956_),
    .B2(\as2650.stack[5][13] ),
    .ZN(_02141_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07766_ (.A1(_02086_),
    .A2(_02140_),
    .A3(_02141_),
    .ZN(_02142_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07767_ (.A1(_02139_),
    .A2(_02142_),
    .B(_01945_),
    .ZN(_02143_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _07768_ (.A1(_02040_),
    .A2(_02135_),
    .B(_02143_),
    .ZN(_02144_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07769_ (.A1(_01934_),
    .A2(_02144_),
    .ZN(_02145_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07770_ (.I(_01533_),
    .Z(_02146_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07771_ (.A1(_02146_),
    .A2(_02099_),
    .ZN(_02147_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _07772_ (.A1(_02071_),
    .A2(_02145_),
    .A3(_02147_),
    .B1(_02101_),
    .B2(_01545_),
    .ZN(_02148_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07773_ (.I0(\as2650.r123[0][5] ),
    .I1(_02148_),
    .S(_02123_),
    .Z(_02149_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07774_ (.I(_02149_),
    .Z(_00035_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07775_ (.A1(\as2650.stack[8][14] ),
    .A2(_02054_),
    .B1(_02037_),
    .B2(\as2650.stack[9][14] ),
    .ZN(_02150_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07776_ (.A1(\as2650.stack[11][14] ),
    .A2(_02029_),
    .B1(_02056_),
    .B2(\as2650.stack[10][14] ),
    .ZN(_02151_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07777_ (.A1(_02079_),
    .A2(_02150_),
    .A3(_02151_),
    .ZN(_02152_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07778_ (.A1(\as2650.stack[15][14] ),
    .A2(_02029_),
    .B1(_02056_),
    .B2(\as2650.stack[14][14] ),
    .ZN(_02153_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07779_ (.A1(\as2650.stack[12][14] ),
    .A2(_02054_),
    .B1(_02037_),
    .B2(\as2650.stack[13][14] ),
    .ZN(_02154_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07780_ (.A1(_02028_),
    .A2(_02153_),
    .A3(_02154_),
    .ZN(_02155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07781_ (.A1(_02152_),
    .A2(_02155_),
    .ZN(_02156_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07782_ (.A1(\as2650.stack[0][14] ),
    .A2(_01814_),
    .B1(_02080_),
    .B2(\as2650.stack[1][14] ),
    .ZN(_02157_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07783_ (.A1(\as2650.stack[3][14] ),
    .A2(_02082_),
    .B1(_02083_),
    .B2(\as2650.stack[2][14] ),
    .ZN(_02158_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07784_ (.A1(_02079_),
    .A2(_02157_),
    .A3(_02158_),
    .ZN(_02159_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07785_ (.A1(\as2650.stack[7][14] ),
    .A2(_02087_),
    .B1(_02126_),
    .B2(\as2650.stack[6][14] ),
    .ZN(_02160_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07786_ (.A1(\as2650.stack[4][14] ),
    .A2(_02089_),
    .B1(_02090_),
    .B2(\as2650.stack[5][14] ),
    .ZN(_02161_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _07787_ (.A1(_02086_),
    .A2(_02160_),
    .A3(_02161_),
    .ZN(_02162_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _07788_ (.A1(_02159_),
    .A2(_02162_),
    .B(_02093_),
    .ZN(_02163_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _07789_ (.A1(_02040_),
    .A2(_02156_),
    .B(_02163_),
    .ZN(_02164_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07790_ (.A1(_01934_),
    .A2(_02164_),
    .ZN(_02165_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07791_ (.A1(_01616_),
    .A2(_02099_),
    .ZN(_02166_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _07792_ (.A1(_02071_),
    .A2(_02165_),
    .A3(_02166_),
    .B1(_02101_),
    .B2(_01636_),
    .ZN(_02167_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07793_ (.I0(\as2650.r123[0][6] ),
    .I1(_02167_),
    .S(_02123_),
    .Z(_02168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07794_ (.I(_02168_),
    .Z(_00036_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _07795_ (.A1(_01921_),
    .A2(_01933_),
    .A3(_01993_),
    .B1(_01718_),
    .B2(_01996_),
    .ZN(_02169_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _07796_ (.I0(\as2650.r123[0][7] ),
    .I1(_02169_),
    .S(_02123_),
    .Z(_02170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07797_ (.I(_02170_),
    .Z(_00037_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07798_ (.I(_01820_),
    .Z(_02171_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07799_ (.I(_01808_),
    .Z(_02172_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07800_ (.I(_01770_),
    .Z(_02173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _07801_ (.A1(_02172_),
    .A2(_02173_),
    .ZN(_02174_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07802_ (.I(_02174_),
    .Z(_02175_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _07803_ (.A1(_01779_),
    .A2(_02171_),
    .A3(_02175_),
    .ZN(_02176_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07804_ (.I(_02176_),
    .Z(_02177_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07805_ (.I(_02177_),
    .Z(_02178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07806_ (.I(_01788_),
    .Z(_02179_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07807_ (.I(_02179_),
    .Z(_02180_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07808_ (.I(_01832_),
    .Z(_02181_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07809_ (.I(net64),
    .Z(_02182_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07810_ (.I(_02182_),
    .Z(_02183_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07811_ (.I(_02183_),
    .Z(_02184_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07812_ (.I(_02184_),
    .Z(_02185_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _07813_ (.A1(_01146_),
    .A2(_02180_),
    .B1(_02181_),
    .B2(_02185_),
    .ZN(_02186_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07814_ (.I(_02186_),
    .Z(_02187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07815_ (.I(_02176_),
    .Z(_02188_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07816_ (.A1(\as2650.stack[14][8] ),
    .A2(_02188_),
    .ZN(_02189_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07817_ (.I(_01766_),
    .Z(_02190_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07818_ (.I(_01824_),
    .Z(_02191_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07819_ (.A1(_02190_),
    .A2(_01778_),
    .A3(_02191_),
    .ZN(_02192_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07820_ (.I(_02192_),
    .Z(_02193_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07821_ (.I(_02193_),
    .Z(_02194_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07822_ (.A1(_02178_),
    .A2(_02187_),
    .B(_02189_),
    .C(_02194_),
    .ZN(_00038_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07823_ (.I(net92),
    .Z(_02195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07824_ (.I(_02195_),
    .Z(_02196_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07825_ (.I(_02196_),
    .Z(_02197_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _07826_ (.A1(_01237_),
    .A2(_02180_),
    .B1(_02181_),
    .B2(_02197_),
    .ZN(_02198_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07827_ (.I(_02198_),
    .Z(_02199_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07828_ (.I(_02176_),
    .Z(_02200_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07829_ (.A1(\as2650.stack[14][9] ),
    .A2(_02200_),
    .ZN(_02201_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07830_ (.A1(_02178_),
    .A2(_02199_),
    .B(_02201_),
    .C(_02194_),
    .ZN(_00039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07831_ (.I(net66),
    .Z(_02202_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07832_ (.I(_02202_),
    .Z(_02203_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07833_ (.I(_02203_),
    .Z(_02204_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _07834_ (.A1(_01313_),
    .A2(_02180_),
    .B1(_02181_),
    .B2(_02204_),
    .ZN(_02205_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07835_ (.I(_02205_),
    .Z(_02206_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07836_ (.A1(\as2650.stack[14][10] ),
    .A2(_02200_),
    .ZN(_02207_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07837_ (.A1(_02178_),
    .A2(_02206_),
    .B(_02207_),
    .C(_02194_),
    .ZN(_00040_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07838_ (.I(net91),
    .Z(_02208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07839_ (.I(_02208_),
    .Z(_02209_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07840_ (.I(_02209_),
    .Z(_02210_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _07841_ (.A1(_01391_),
    .A2(_02180_),
    .B1(_02181_),
    .B2(_02210_),
    .ZN(_02211_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07842_ (.I(_02211_),
    .Z(_02212_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07843_ (.A1(\as2650.stack[14][11] ),
    .A2(_02200_),
    .ZN(_02213_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07844_ (.A1(_02178_),
    .A2(_02212_),
    .B(_02213_),
    .C(_02194_),
    .ZN(_00041_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07845_ (.I(_02177_),
    .Z(_02214_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07846_ (.I(net68),
    .Z(_02215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07847_ (.I(_02215_),
    .Z(_02216_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07848_ (.I(_02216_),
    .Z(_02217_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _07849_ (.A1(_01724_),
    .A2(_02179_),
    .B1(_01833_),
    .B2(_02217_),
    .ZN(_02218_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07850_ (.I(_02218_),
    .Z(_02219_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07851_ (.A1(\as2650.stack[14][12] ),
    .A2(_02200_),
    .ZN(_02220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07852_ (.I(_02193_),
    .Z(_02221_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07853_ (.A1(_02214_),
    .A2(_02219_),
    .B(_02220_),
    .C(_02221_),
    .ZN(_00042_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07854_ (.I(_01733_),
    .Z(_02222_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07855_ (.I(_02222_),
    .Z(_02223_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07856_ (.I(net69),
    .Z(_02224_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _07857_ (.A1(_02223_),
    .A2(_02179_),
    .B1(_01833_),
    .B2(_02224_),
    .ZN(_02225_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07858_ (.I(_02225_),
    .Z(_02226_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07859_ (.A1(\as2650.stack[14][13] ),
    .A2(_02177_),
    .ZN(_02227_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07860_ (.A1(_02214_),
    .A2(_02226_),
    .B(_02227_),
    .C(_02221_),
    .ZN(_00043_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07861_ (.I(_01742_),
    .Z(_02228_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07862_ (.I(_02228_),
    .Z(_02229_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07863_ (.I(_02229_),
    .Z(_02230_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _07864_ (.I(net71),
    .Z(_02231_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _07865_ (.A1(_02230_),
    .A2(_02179_),
    .B1(_01833_),
    .B2(_02231_),
    .ZN(_02232_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07866_ (.I(_02232_),
    .Z(_02233_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07867_ (.A1(\as2650.stack[14][14] ),
    .A2(_02177_),
    .ZN(_02234_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07868_ (.A1(_02214_),
    .A2(_02233_),
    .B(_02234_),
    .C(_02221_),
    .ZN(_00044_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07869_ (.I(_01827_),
    .Z(_02235_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07870_ (.A1(\as2650.stack[13][8] ),
    .A2(_01898_),
    .ZN(_02236_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07871_ (.I(_01841_),
    .Z(_02237_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07872_ (.A1(_02235_),
    .A2(_02187_),
    .B(_02236_),
    .C(_02237_),
    .ZN(_00045_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07873_ (.I(_01826_),
    .Z(_02238_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07874_ (.A1(\as2650.stack[13][9] ),
    .A2(_02238_),
    .ZN(_02239_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07875_ (.A1(_02235_),
    .A2(_02199_),
    .B(_02239_),
    .C(_02237_),
    .ZN(_00046_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07876_ (.A1(\as2650.stack[13][10] ),
    .A2(_02238_),
    .ZN(_02240_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07877_ (.A1(_02235_),
    .A2(_02206_),
    .B(_02240_),
    .C(_02237_),
    .ZN(_00047_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07878_ (.A1(\as2650.stack[13][11] ),
    .A2(_02238_),
    .ZN(_02241_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07879_ (.A1(_02235_),
    .A2(_02212_),
    .B(_02241_),
    .C(_02237_),
    .ZN(_00048_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07880_ (.A1(\as2650.stack[13][12] ),
    .A2(_02238_),
    .ZN(_02242_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07881_ (.A1(_01828_),
    .A2(_02219_),
    .B(_02242_),
    .C(_01842_),
    .ZN(_00049_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07882_ (.A1(\as2650.stack[13][13] ),
    .A2(_01827_),
    .ZN(_02243_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07883_ (.A1(_01828_),
    .A2(_02226_),
    .B(_02243_),
    .C(_01842_),
    .ZN(_00050_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07884_ (.A1(\as2650.stack[13][14] ),
    .A2(_01827_),
    .ZN(_02244_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07885_ (.A1(_01828_),
    .A2(_02233_),
    .B(_02244_),
    .C(_01842_),
    .ZN(_00051_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07886_ (.I(_01937_),
    .Z(_02245_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07887_ (.I(_02245_),
    .Z(_02246_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07888_ (.A1(_02190_),
    .A2(_02191_),
    .A3(_02246_),
    .ZN(_02247_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07889_ (.I(_02247_),
    .Z(_02248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07890_ (.I(_02248_),
    .Z(_02249_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07891_ (.I(_01806_),
    .Z(_02250_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _07892_ (.I(_01776_),
    .ZN(_02251_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07893_ (.A1(_01774_),
    .A2(_02251_),
    .ZN(_02252_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07894_ (.I(_02252_),
    .Z(_02253_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07895_ (.I(_02080_),
    .Z(_02254_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07896_ (.I(_02254_),
    .Z(_02255_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _07897_ (.A1(_02250_),
    .A2(_02253_),
    .A3(_02255_),
    .ZN(_02256_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07898_ (.I(_02256_),
    .Z(_02257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07899_ (.A1(\as2650.stack[10][0] ),
    .A2(_02257_),
    .ZN(_02258_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _07900_ (.I(_01839_),
    .Z(_02259_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07901_ (.I(_02171_),
    .Z(_02260_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _07902_ (.A1(_02260_),
    .A2(_02246_),
    .A3(_02175_),
    .ZN(_02261_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07903_ (.I(_02261_),
    .Z(_02262_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07904_ (.I(_02262_),
    .Z(_02263_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07905_ (.I(_02247_),
    .Z(_02264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07906_ (.I(_02264_),
    .Z(_02265_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _07907_ (.A1(_02259_),
    .A2(_02263_),
    .B(_02265_),
    .ZN(_02266_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07908_ (.A1(_01762_),
    .A2(_02249_),
    .B1(_02258_),
    .B2(_02266_),
    .ZN(_00052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07909_ (.A1(\as2650.stack[10][1] ),
    .A2(_02257_),
    .ZN(_02267_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07910_ (.I(_01857_),
    .Z(_02268_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07911_ (.I(_02261_),
    .Z(_02269_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07912_ (.I(_02264_),
    .Z(_02270_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07913_ (.A1(_02268_),
    .A2(_02269_),
    .B(_02270_),
    .ZN(_02271_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07914_ (.A1(_01847_),
    .A2(_02249_),
    .B1(_02267_),
    .B2(_02271_),
    .ZN(_00053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07915_ (.A1(\as2650.stack[10][2] ),
    .A2(_02257_),
    .ZN(_02272_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07916_ (.I(_01869_),
    .Z(_02273_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07917_ (.A1(_02273_),
    .A2(_02269_),
    .B(_02270_),
    .ZN(_02274_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07918_ (.A1(_01863_),
    .A2(_02249_),
    .B1(_02272_),
    .B2(_02274_),
    .ZN(_00054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07919_ (.A1(\as2650.stack[10][3] ),
    .A2(_02257_),
    .ZN(_02275_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07920_ (.I(_01880_),
    .Z(_02276_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07921_ (.A1(_02276_),
    .A2(_02269_),
    .B(_02270_),
    .ZN(_02277_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07922_ (.A1(_01874_),
    .A2(_02249_),
    .B1(_02275_),
    .B2(_02277_),
    .ZN(_00055_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07923_ (.I(_02264_),
    .Z(_02278_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07924_ (.I(_02256_),
    .Z(_02279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07925_ (.A1(\as2650.stack[10][4] ),
    .A2(_02279_),
    .ZN(_02280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07926_ (.I(_01891_),
    .Z(_02281_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07927_ (.A1(_02281_),
    .A2(_02269_),
    .B(_02270_),
    .ZN(_02282_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07928_ (.A1(_01884_),
    .A2(_02278_),
    .B1(_02280_),
    .B2(_02282_),
    .ZN(_00056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07929_ (.A1(\as2650.stack[10][5] ),
    .A2(_02279_),
    .ZN(_02283_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07930_ (.I(_01905_),
    .Z(_02284_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07931_ (.I(_02261_),
    .Z(_02285_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07932_ (.A1(_02284_),
    .A2(_02285_),
    .B(_02248_),
    .ZN(_02286_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07933_ (.A1(_01896_),
    .A2(_02278_),
    .B1(_02283_),
    .B2(_02286_),
    .ZN(_00057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07934_ (.A1(\as2650.stack[10][6] ),
    .A2(_02279_),
    .ZN(_02287_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07935_ (.I(_01915_),
    .Z(_02288_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07936_ (.A1(_02288_),
    .A2(_02285_),
    .B(_02248_),
    .ZN(_02289_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07937_ (.A1(_01909_),
    .A2(_02278_),
    .B1(_02287_),
    .B2(_02289_),
    .ZN(_00058_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07938_ (.A1(\as2650.stack[10][7] ),
    .A2(_02279_),
    .ZN(_02290_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07939_ (.I(_01924_),
    .Z(_02291_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _07940_ (.A1(_02291_),
    .A2(_02285_),
    .B(_02248_),
    .ZN(_02292_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _07941_ (.A1(_01919_),
    .A2(_02278_),
    .B1(_02290_),
    .B2(_02292_),
    .ZN(_00059_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _07942_ (.A1(_01772_),
    .A2(_01779_),
    .A3(_02260_),
    .ZN(_02293_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07943_ (.I(_02293_),
    .Z(_02294_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07944_ (.I(_02294_),
    .Z(_02295_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07945_ (.I(_02293_),
    .Z(_02296_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07946_ (.A1(\as2650.stack[12][8] ),
    .A2(_02296_),
    .ZN(_02297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _07947_ (.A1(_01808_),
    .A2(_01823_),
    .ZN(_02298_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07948_ (.I(_02298_),
    .Z(_02299_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _07949_ (.A1(_02190_),
    .A2(_02245_),
    .A3(_02299_),
    .ZN(_02300_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07950_ (.I(_02300_),
    .Z(_02301_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07951_ (.I(_02301_),
    .Z(_02302_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07952_ (.A1(_02187_),
    .A2(_02295_),
    .B(_02297_),
    .C(_02302_),
    .ZN(_00060_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07953_ (.I(_02293_),
    .Z(_02303_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07954_ (.A1(\as2650.stack[12][9] ),
    .A2(_02303_),
    .ZN(_02304_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07955_ (.A1(_02199_),
    .A2(_02295_),
    .B(_02304_),
    .C(_02302_),
    .ZN(_00061_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07956_ (.A1(\as2650.stack[12][10] ),
    .A2(_02303_),
    .ZN(_02305_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07957_ (.A1(_02206_),
    .A2(_02295_),
    .B(_02305_),
    .C(_02302_),
    .ZN(_00062_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07958_ (.A1(\as2650.stack[12][11] ),
    .A2(_02303_),
    .ZN(_02306_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07959_ (.A1(_02212_),
    .A2(_02295_),
    .B(_02306_),
    .C(_02302_),
    .ZN(_00063_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07960_ (.I(_02294_),
    .Z(_02307_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07961_ (.A1(\as2650.stack[12][12] ),
    .A2(_02303_),
    .ZN(_02308_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07962_ (.I(_02301_),
    .Z(_02309_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07963_ (.A1(_02219_),
    .A2(_02307_),
    .B(_02308_),
    .C(_02309_),
    .ZN(_00064_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07964_ (.A1(\as2650.stack[12][13] ),
    .A2(_02294_),
    .ZN(_02310_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07965_ (.A1(_02226_),
    .A2(_02307_),
    .B(_02310_),
    .C(_02309_),
    .ZN(_00065_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07966_ (.A1(\as2650.stack[12][14] ),
    .A2(_02294_),
    .ZN(_02311_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07967_ (.A1(_02233_),
    .A2(_02307_),
    .B(_02311_),
    .C(_02309_),
    .ZN(_00066_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _07968_ (.I(_02171_),
    .Z(_02312_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _07969_ (.A1(_02312_),
    .A2(_02246_),
    .A3(_02299_),
    .ZN(_02313_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07970_ (.I(_02313_),
    .Z(_02314_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07971_ (.I(_02314_),
    .Z(_02315_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07972_ (.I(_02313_),
    .Z(_02316_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07973_ (.A1(\as2650.stack[11][8] ),
    .A2(_02316_),
    .ZN(_02317_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07974_ (.I(_02174_),
    .Z(_02318_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _07975_ (.A1(_02190_),
    .A2(_02245_),
    .A3(_02318_),
    .ZN(_02319_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07976_ (.I(_02319_),
    .Z(_02320_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07977_ (.I(_02320_),
    .Z(_02321_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07978_ (.A1(_02187_),
    .A2(_02315_),
    .B(_02317_),
    .C(_02321_),
    .ZN(_00067_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07979_ (.I(_02313_),
    .Z(_02322_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07980_ (.A1(\as2650.stack[11][9] ),
    .A2(_02322_),
    .ZN(_02323_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07981_ (.A1(_02199_),
    .A2(_02315_),
    .B(_02323_),
    .C(_02321_),
    .ZN(_00068_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07982_ (.A1(\as2650.stack[11][10] ),
    .A2(_02322_),
    .ZN(_02324_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07983_ (.A1(_02206_),
    .A2(_02315_),
    .B(_02324_),
    .C(_02321_),
    .ZN(_00069_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07984_ (.A1(\as2650.stack[11][11] ),
    .A2(_02322_),
    .ZN(_02325_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07985_ (.A1(_02212_),
    .A2(_02315_),
    .B(_02325_),
    .C(_02321_),
    .ZN(_00070_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _07986_ (.I(_02314_),
    .Z(_02326_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07987_ (.A1(\as2650.stack[11][12] ),
    .A2(_02322_),
    .ZN(_02327_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _07988_ (.I(_02320_),
    .Z(_02328_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07989_ (.A1(_02219_),
    .A2(_02326_),
    .B(_02327_),
    .C(_02328_),
    .ZN(_00071_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07990_ (.A1(\as2650.stack[11][13] ),
    .A2(_02314_),
    .ZN(_02329_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07991_ (.A1(_02226_),
    .A2(_02326_),
    .B(_02329_),
    .C(_02328_),
    .ZN(_00072_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07992_ (.A1(\as2650.stack[11][14] ),
    .A2(_02314_),
    .ZN(_02330_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _07993_ (.A1(_02233_),
    .A2(_02326_),
    .B(_02330_),
    .C(_02328_),
    .ZN(_00073_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _07994_ (.A1(_00779_),
    .A2(_00574_),
    .ZN(_02331_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _07995_ (.I(_02331_),
    .ZN(_02332_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _07996_ (.A1(_00836_),
    .A2(_02332_),
    .ZN(_02333_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _07997_ (.I(_01793_),
    .Z(_02334_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _07998_ (.I(_02334_),
    .Z(_02335_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _07999_ (.A1(_00500_),
    .A2(_00567_),
    .ZN(_02336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08000_ (.A1(_00509_),
    .A2(_00874_),
    .ZN(_02337_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08001_ (.A1(_00971_),
    .A2(_02337_),
    .ZN(_02338_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08002_ (.A1(_02336_),
    .A2(_02338_),
    .Z(_02339_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08003_ (.I(_02339_),
    .Z(_02340_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08004_ (.A1(_00584_),
    .A2(_00944_),
    .B1(_02335_),
    .B2(_02340_),
    .ZN(_02341_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08005_ (.I(_02341_),
    .ZN(_02342_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08006_ (.A1(_02333_),
    .A2(_02342_),
    .ZN(_02343_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08007_ (.A1(_00936_),
    .A2(_00948_),
    .A3(_00949_),
    .ZN(_02344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08008_ (.A1(_01703_),
    .A2(_00535_),
    .ZN(_02345_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08009_ (.I(net77),
    .ZN(_02346_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08010_ (.I(_00972_),
    .Z(_02347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08011_ (.A1(_02347_),
    .A2(_00851_),
    .ZN(_02348_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08012_ (.A1(_00851_),
    .A2(_02346_),
    .B(_02348_),
    .ZN(_02349_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08013_ (.A1(_02335_),
    .A2(_02340_),
    .A3(_02349_),
    .ZN(_02350_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08014_ (.A1(_02344_),
    .A2(_02345_),
    .B(_02350_),
    .ZN(_02351_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08015_ (.A1(net4),
    .A2(_02343_),
    .B1(_02351_),
    .B2(_02333_),
    .ZN(_02352_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08016_ (.A1(_00773_),
    .A2(_02352_),
    .ZN(_00074_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08017_ (.I(_02192_),
    .Z(_02353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08018_ (.I(_02353_),
    .Z(_02354_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _08019_ (.A1(_01783_),
    .A2(_01785_),
    .A3(_01807_),
    .A4(_02255_),
    .ZN(_02355_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08020_ (.I(_02355_),
    .Z(_02356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08021_ (.A1(\as2650.stack[14][0] ),
    .A2(_02356_),
    .ZN(_02357_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08022_ (.A1(_02259_),
    .A2(_02214_),
    .B(_02221_),
    .ZN(_02358_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08023_ (.A1(_01762_),
    .A2(_02354_),
    .B1(_02357_),
    .B2(_02358_),
    .ZN(_00075_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08024_ (.A1(\as2650.stack[14][1] ),
    .A2(_02356_),
    .ZN(_02359_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08025_ (.I(_02176_),
    .Z(_02360_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08026_ (.I(_02193_),
    .Z(_02361_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08027_ (.A1(_02268_),
    .A2(_02360_),
    .B(_02361_),
    .ZN(_02362_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08028_ (.A1(_01847_),
    .A2(_02354_),
    .B1(_02359_),
    .B2(_02362_),
    .ZN(_00076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08029_ (.A1(\as2650.stack[14][2] ),
    .A2(_02356_),
    .ZN(_02363_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08030_ (.A1(_02273_),
    .A2(_02360_),
    .B(_02361_),
    .ZN(_02364_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08031_ (.A1(_01863_),
    .A2(_02354_),
    .B1(_02363_),
    .B2(_02364_),
    .ZN(_00077_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08032_ (.A1(\as2650.stack[14][3] ),
    .A2(_02356_),
    .ZN(_02365_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08033_ (.A1(_02276_),
    .A2(_02360_),
    .B(_02361_),
    .ZN(_02366_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08034_ (.A1(_01874_),
    .A2(_02354_),
    .B1(_02365_),
    .B2(_02366_),
    .ZN(_00078_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08035_ (.I(_02193_),
    .Z(_02367_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08036_ (.I(_02355_),
    .Z(_02368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08037_ (.A1(\as2650.stack[14][4] ),
    .A2(_02368_),
    .ZN(_02369_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08038_ (.A1(_02281_),
    .A2(_02360_),
    .B(_02361_),
    .ZN(_02370_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08039_ (.A1(_01884_),
    .A2(_02367_),
    .B1(_02369_),
    .B2(_02370_),
    .ZN(_00079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08040_ (.A1(\as2650.stack[14][5] ),
    .A2(_02368_),
    .ZN(_02371_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08041_ (.A1(_02284_),
    .A2(_02188_),
    .B(_02353_),
    .ZN(_02372_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08042_ (.A1(_01896_),
    .A2(_02367_),
    .B1(_02371_),
    .B2(_02372_),
    .ZN(_00080_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08043_ (.A1(\as2650.stack[14][6] ),
    .A2(_02368_),
    .ZN(_02373_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08044_ (.A1(_02288_),
    .A2(_02188_),
    .B(_02353_),
    .ZN(_02374_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08045_ (.A1(_01909_),
    .A2(_02367_),
    .B1(_02373_),
    .B2(_02374_),
    .ZN(_00081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08046_ (.A1(\as2650.stack[14][7] ),
    .A2(_02368_),
    .ZN(_02375_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08047_ (.A1(_02291_),
    .A2(_02188_),
    .B(_02353_),
    .ZN(_02376_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08048_ (.A1(_01919_),
    .A2(_02367_),
    .B1(_02375_),
    .B2(_02376_),
    .ZN(_00082_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08049_ (.I(_02186_),
    .Z(_02377_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08050_ (.I(_02262_),
    .Z(_02378_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08051_ (.A1(\as2650.stack[10][8] ),
    .A2(_02285_),
    .ZN(_02379_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08052_ (.I(_02264_),
    .Z(_02380_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08053_ (.A1(_02377_),
    .A2(_02378_),
    .B(_02379_),
    .C(_02380_),
    .ZN(_00083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08054_ (.I(_02198_),
    .Z(_02381_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08055_ (.I(_02261_),
    .Z(_02382_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08056_ (.A1(\as2650.stack[10][9] ),
    .A2(_02382_),
    .ZN(_02383_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08057_ (.A1(_02381_),
    .A2(_02378_),
    .B(_02383_),
    .C(_02380_),
    .ZN(_00084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08058_ (.I(_02205_),
    .Z(_02384_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08059_ (.A1(\as2650.stack[10][10] ),
    .A2(_02382_),
    .ZN(_02385_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08060_ (.A1(_02384_),
    .A2(_02378_),
    .B(_02385_),
    .C(_02380_),
    .ZN(_00085_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08061_ (.I(_02211_),
    .Z(_02386_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08062_ (.A1(\as2650.stack[10][11] ),
    .A2(_02382_),
    .ZN(_02387_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08063_ (.A1(_02386_),
    .A2(_02378_),
    .B(_02387_),
    .C(_02380_),
    .ZN(_00086_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08064_ (.I(_02218_),
    .Z(_02388_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08065_ (.A1(\as2650.stack[10][12] ),
    .A2(_02382_),
    .ZN(_02389_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08066_ (.A1(_02388_),
    .A2(_02263_),
    .B(_02389_),
    .C(_02265_),
    .ZN(_00087_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08067_ (.I(_02225_),
    .Z(_02390_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08068_ (.A1(\as2650.stack[10][13] ),
    .A2(_02262_),
    .ZN(_02391_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08069_ (.A1(_02390_),
    .A2(_02263_),
    .B(_02391_),
    .C(_02265_),
    .ZN(_00088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08070_ (.I(_02232_),
    .Z(_02392_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08071_ (.A1(\as2650.stack[10][14] ),
    .A2(_02262_),
    .ZN(_02393_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08072_ (.A1(_02392_),
    .A2(_02263_),
    .B(_02393_),
    .C(_02265_),
    .ZN(_00089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08073_ (.I(_02137_),
    .Z(_02394_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08074_ (.A1(_01783_),
    .A2(_01784_),
    .A3(_02394_),
    .ZN(_02395_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08075_ (.A1(_01767_),
    .A2(_02395_),
    .ZN(_02396_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08076_ (.I(_02396_),
    .Z(_02397_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08077_ (.I(_02397_),
    .Z(_02398_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08078_ (.I(_02007_),
    .Z(_02399_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08079_ (.I(_01806_),
    .Z(_02400_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08080_ (.A1(_01775_),
    .A2(_01784_),
    .ZN(_02401_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08081_ (.I(_02401_),
    .Z(_02402_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _08082_ (.A1(_02399_),
    .A2(_02400_),
    .A3(_02402_),
    .ZN(_02403_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08083_ (.I(_02403_),
    .Z(_02404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08084_ (.A1(\as2650.stack[0][0] ),
    .A2(_02404_),
    .ZN(_02405_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08085_ (.I(_01936_),
    .Z(_02406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08086_ (.A1(_02406_),
    .A2(_02251_),
    .ZN(_02407_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08087_ (.I(_02407_),
    .Z(_02408_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _08088_ (.A1(_01772_),
    .A2(_02260_),
    .A3(_02408_),
    .ZN(_02409_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08089_ (.I(_02409_),
    .Z(_02410_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08090_ (.I(_02410_),
    .Z(_02411_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08091_ (.I(_02396_),
    .Z(_02412_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08092_ (.I(_02412_),
    .Z(_02413_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08093_ (.A1(_02259_),
    .A2(_02411_),
    .B(_02413_),
    .ZN(_02414_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08094_ (.A1(_01762_),
    .A2(_02398_),
    .B1(_02405_),
    .B2(_02414_),
    .ZN(_00090_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08095_ (.A1(\as2650.stack[0][1] ),
    .A2(_02404_),
    .ZN(_02415_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08096_ (.I(_02409_),
    .Z(_02416_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08097_ (.I(_02412_),
    .Z(_02417_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08098_ (.A1(_02268_),
    .A2(_02416_),
    .B(_02417_),
    .ZN(_02418_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08099_ (.A1(_01847_),
    .A2(_02398_),
    .B1(_02415_),
    .B2(_02418_),
    .ZN(_00091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08100_ (.A1(\as2650.stack[0][2] ),
    .A2(_02404_),
    .ZN(_02419_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08101_ (.A1(_02273_),
    .A2(_02416_),
    .B(_02417_),
    .ZN(_02420_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08102_ (.A1(_01863_),
    .A2(_02398_),
    .B1(_02419_),
    .B2(_02420_),
    .ZN(_00092_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08103_ (.A1(\as2650.stack[0][3] ),
    .A2(_02404_),
    .ZN(_02421_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08104_ (.A1(_02276_),
    .A2(_02416_),
    .B(_02417_),
    .ZN(_02422_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08105_ (.A1(_01874_),
    .A2(_02398_),
    .B1(_02421_),
    .B2(_02422_),
    .ZN(_00093_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08106_ (.I(_02412_),
    .Z(_02423_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08107_ (.I(_02403_),
    .Z(_02424_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08108_ (.A1(\as2650.stack[0][4] ),
    .A2(_02424_),
    .ZN(_02425_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08109_ (.A1(_02281_),
    .A2(_02416_),
    .B(_02417_),
    .ZN(_02426_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08110_ (.A1(_01884_),
    .A2(_02423_),
    .B1(_02425_),
    .B2(_02426_),
    .ZN(_00094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08111_ (.A1(\as2650.stack[0][5] ),
    .A2(_02424_),
    .ZN(_02427_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08112_ (.I(_02409_),
    .Z(_02428_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08113_ (.A1(_02284_),
    .A2(_02428_),
    .B(_02397_),
    .ZN(_02429_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08114_ (.A1(_01896_),
    .A2(_02423_),
    .B1(_02427_),
    .B2(_02429_),
    .ZN(_00095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08115_ (.A1(\as2650.stack[0][6] ),
    .A2(_02424_),
    .ZN(_02430_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08116_ (.A1(_02288_),
    .A2(_02428_),
    .B(_02397_),
    .ZN(_02431_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08117_ (.A1(_01909_),
    .A2(_02423_),
    .B1(_02430_),
    .B2(_02431_),
    .ZN(_00096_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08118_ (.A1(\as2650.stack[0][7] ),
    .A2(_02424_),
    .ZN(_02432_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08119_ (.A1(_02291_),
    .A2(_02428_),
    .B(_02397_),
    .ZN(_02433_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08120_ (.A1(_01919_),
    .A2(_02423_),
    .B1(_02432_),
    .B2(_02433_),
    .ZN(_00097_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08121_ (.I(_02410_),
    .Z(_02434_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08122_ (.A1(\as2650.stack[0][8] ),
    .A2(_02428_),
    .ZN(_02435_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08123_ (.I(_02412_),
    .Z(_02436_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08124_ (.A1(_02377_),
    .A2(_02434_),
    .B(_02435_),
    .C(_02436_),
    .ZN(_00098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08125_ (.I(_02409_),
    .Z(_02437_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08126_ (.A1(\as2650.stack[0][9] ),
    .A2(_02437_),
    .ZN(_02438_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08127_ (.A1(_02381_),
    .A2(_02434_),
    .B(_02438_),
    .C(_02436_),
    .ZN(_00099_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08128_ (.A1(\as2650.stack[0][10] ),
    .A2(_02437_),
    .ZN(_02439_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08129_ (.A1(_02384_),
    .A2(_02434_),
    .B(_02439_),
    .C(_02436_),
    .ZN(_00100_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08130_ (.A1(\as2650.stack[0][11] ),
    .A2(_02437_),
    .ZN(_02440_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08131_ (.A1(_02386_),
    .A2(_02434_),
    .B(_02440_),
    .C(_02436_),
    .ZN(_00101_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08132_ (.A1(\as2650.stack[0][12] ),
    .A2(_02437_),
    .ZN(_02441_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08133_ (.A1(_02388_),
    .A2(_02411_),
    .B(_02441_),
    .C(_02413_),
    .ZN(_00102_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08134_ (.A1(\as2650.stack[0][13] ),
    .A2(_02410_),
    .ZN(_02442_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08135_ (.A1(_02390_),
    .A2(_02411_),
    .B(_02442_),
    .C(_02413_),
    .ZN(_00103_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08136_ (.A1(\as2650.stack[0][14] ),
    .A2(_02410_),
    .ZN(_02443_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08137_ (.A1(_02392_),
    .A2(_02411_),
    .B(_02443_),
    .C(_02413_),
    .ZN(_00104_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08138_ (.I(_02171_),
    .Z(_02444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08139_ (.A1(_02007_),
    .A2(_02253_),
    .ZN(_02445_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08140_ (.A1(_02444_),
    .A2(_02445_),
    .ZN(_02446_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08141_ (.I(_02446_),
    .Z(_02447_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08142_ (.I(_02447_),
    .Z(_02448_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08143_ (.I(_02446_),
    .Z(_02449_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08144_ (.A1(\as2650.stack[8][8] ),
    .A2(_02449_),
    .ZN(_02450_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08145_ (.I(_01766_),
    .Z(_02451_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08146_ (.A1(_01775_),
    .A2(_02251_),
    .ZN(_02452_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08147_ (.I(_02452_),
    .Z(_02453_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08148_ (.A1(_02451_),
    .A2(_02299_),
    .A3(_02453_),
    .ZN(_02454_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08149_ (.I(_02454_),
    .Z(_02455_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08150_ (.I(_02455_),
    .Z(_02456_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08151_ (.A1(_02377_),
    .A2(_02448_),
    .B(_02450_),
    .C(_02456_),
    .ZN(_00105_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08152_ (.I(_02446_),
    .Z(_02457_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08153_ (.A1(\as2650.stack[8][9] ),
    .A2(_02457_),
    .ZN(_02458_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08154_ (.A1(_02381_),
    .A2(_02448_),
    .B(_02458_),
    .C(_02456_),
    .ZN(_00106_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08155_ (.A1(\as2650.stack[8][10] ),
    .A2(_02457_),
    .ZN(_02459_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08156_ (.A1(_02384_),
    .A2(_02448_),
    .B(_02459_),
    .C(_02456_),
    .ZN(_00107_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08157_ (.A1(\as2650.stack[8][11] ),
    .A2(_02457_),
    .ZN(_02460_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08158_ (.A1(_02386_),
    .A2(_02448_),
    .B(_02460_),
    .C(_02456_),
    .ZN(_00108_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08159_ (.I(_02447_),
    .Z(_02461_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08160_ (.A1(\as2650.stack[8][12] ),
    .A2(_02457_),
    .ZN(_02462_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08161_ (.I(_02455_),
    .Z(_02463_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08162_ (.A1(_02388_),
    .A2(_02461_),
    .B(_02462_),
    .C(_02463_),
    .ZN(_00109_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08163_ (.A1(\as2650.stack[8][13] ),
    .A2(_02447_),
    .ZN(_02464_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08164_ (.A1(_02390_),
    .A2(_02461_),
    .B(_02464_),
    .C(_02463_),
    .ZN(_00110_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08165_ (.A1(\as2650.stack[8][14] ),
    .A2(_02447_),
    .ZN(_02465_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08166_ (.A1(_02392_),
    .A2(_02461_),
    .B(_02465_),
    .C(_02463_),
    .ZN(_00111_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08167_ (.I(_02452_),
    .Z(_02466_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _08168_ (.A1(_02312_),
    .A2(_02299_),
    .A3(_02466_),
    .ZN(_02467_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08169_ (.I(_02467_),
    .Z(_02468_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08170_ (.I(_02468_),
    .Z(_02469_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08171_ (.I(_02467_),
    .Z(_02470_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08172_ (.A1(\as2650.stack[7][8] ),
    .A2(_02470_),
    .ZN(_02471_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08173_ (.A1(_02451_),
    .A2(_02318_),
    .A3(_02453_),
    .ZN(_02472_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08174_ (.I(_02472_),
    .Z(_02473_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08175_ (.I(_02473_),
    .Z(_02474_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08176_ (.A1(_02377_),
    .A2(_02469_),
    .B(_02471_),
    .C(_02474_),
    .ZN(_00112_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08177_ (.I(_02467_),
    .Z(_02475_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08178_ (.A1(\as2650.stack[7][9] ),
    .A2(_02475_),
    .ZN(_02476_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08179_ (.A1(_02381_),
    .A2(_02469_),
    .B(_02476_),
    .C(_02474_),
    .ZN(_00113_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08180_ (.A1(\as2650.stack[7][10] ),
    .A2(_02475_),
    .ZN(_02477_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08181_ (.A1(_02384_),
    .A2(_02469_),
    .B(_02477_),
    .C(_02474_),
    .ZN(_00114_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08182_ (.A1(\as2650.stack[7][11] ),
    .A2(_02475_),
    .ZN(_02478_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08183_ (.A1(_02386_),
    .A2(_02469_),
    .B(_02478_),
    .C(_02474_),
    .ZN(_00115_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08184_ (.I(_02468_),
    .Z(_02479_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08185_ (.A1(\as2650.stack[7][12] ),
    .A2(_02475_),
    .ZN(_02480_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08186_ (.I(_02473_),
    .Z(_02481_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08187_ (.A1(_02388_),
    .A2(_02479_),
    .B(_02480_),
    .C(_02481_),
    .ZN(_00116_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08188_ (.A1(\as2650.stack[7][13] ),
    .A2(_02468_),
    .ZN(_02482_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08189_ (.A1(_02390_),
    .A2(_02479_),
    .B(_02482_),
    .C(_02481_),
    .ZN(_00117_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08190_ (.A1(\as2650.stack[7][14] ),
    .A2(_02468_),
    .ZN(_02483_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08191_ (.A1(_02392_),
    .A2(_02479_),
    .B(_02483_),
    .C(_02481_),
    .ZN(_00118_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08192_ (.I(net75),
    .Z(_02484_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08193_ (.I(_02484_),
    .ZN(_02485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08194_ (.I(_00992_),
    .Z(_02486_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08195_ (.A1(_00572_),
    .A2(_01928_),
    .A3(_00981_),
    .A4(_02486_),
    .Z(_02487_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _08196_ (.A1(_02347_),
    .A2(_00949_),
    .A3(_00964_),
    .ZN(_02488_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _08197_ (.A1(_02344_),
    .A2(_00975_),
    .A3(_02487_),
    .A4(_02488_),
    .ZN(_02489_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _08198_ (.A1(_00672_),
    .A2(_00905_),
    .ZN(_02490_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08199_ (.A1(_00832_),
    .A2(_00563_),
    .ZN(_02491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08200_ (.A1(_02490_),
    .A2(_02491_),
    .ZN(_02492_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _08201_ (.A1(_00533_),
    .A2(_02492_),
    .A3(_00571_),
    .A4(_02332_),
    .ZN(_02493_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08202_ (.I(_02336_),
    .Z(_02494_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08203_ (.A1(_00971_),
    .A2(_00482_),
    .ZN(_02495_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08204_ (.A1(_00972_),
    .A2(_02495_),
    .ZN(_02496_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08205_ (.A1(_02494_),
    .A2(_02496_),
    .Z(_02497_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08206_ (.A1(_00582_),
    .A2(_02340_),
    .A3(_02497_),
    .ZN(_02498_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08207_ (.A1(_00899_),
    .A2(_02493_),
    .A3(_02498_),
    .ZN(_02499_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _08208_ (.A1(_00781_),
    .A2(_00725_),
    .ZN(_02500_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08209_ (.A1(_00995_),
    .A2(_02500_),
    .ZN(_02501_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08210_ (.A1(_00780_),
    .A2(_00502_),
    .ZN(_02502_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08211_ (.A1(_00529_),
    .A2(_02500_),
    .B1(_02502_),
    .B2(_00498_),
    .ZN(_02503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _08212_ (.A1(_02501_),
    .A2(_02503_),
    .ZN(_02504_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _08213_ (.A1(_02494_),
    .A2(_02496_),
    .ZN(_02505_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08214_ (.A1(_00717_),
    .A2(_00576_),
    .A3(_00858_),
    .ZN(_02506_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08215_ (.A1(_05721_),
    .A2(_00497_),
    .ZN(_02507_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _08216_ (.A1(_00779_),
    .A2(_00579_),
    .ZN(_02508_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08217_ (.A1(_02507_),
    .A2(_02508_),
    .ZN(_02509_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08218_ (.A1(_02505_),
    .A2(_02506_),
    .A3(_02509_),
    .ZN(_02510_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08219_ (.A1(_02504_),
    .A2(_02510_),
    .ZN(_02511_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08220_ (.A1(_02489_),
    .A2(_02499_),
    .A3(_02511_),
    .ZN(_02512_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08221_ (.I(_00571_),
    .ZN(_02513_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08222_ (.A1(_00579_),
    .A2(_00673_),
    .ZN(_02514_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08223_ (.I(_02514_),
    .Z(_02515_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08224_ (.I(_02515_),
    .Z(_02516_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _08225_ (.A1(_00682_),
    .A2(_02513_),
    .A3(_02516_),
    .A4(_02500_),
    .ZN(_02517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08226_ (.A1(_00563_),
    .A2(_02486_),
    .ZN(_02518_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _08227_ (.A1(_00780_),
    .A2(_00655_),
    .ZN(_02519_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _08228_ (.A1(_05746_),
    .A2(_00954_),
    .A3(_02518_),
    .B1(_02519_),
    .B2(_00966_),
    .ZN(_02520_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08229_ (.A1(_00749_),
    .A2(_00690_),
    .ZN(_02521_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08230_ (.A1(_00832_),
    .A2(_01016_),
    .ZN(_02522_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08231_ (.A1(_01399_),
    .A2(_02522_),
    .A3(_02333_),
    .ZN(_02523_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08232_ (.I(_02523_),
    .ZN(_02524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _08233_ (.A1(_00797_),
    .A2(_00532_),
    .ZN(_02525_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _08234_ (.A1(_01061_),
    .A2(_00934_),
    .A3(_00981_),
    .A4(_02525_),
    .ZN(_02526_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _08235_ (.A1(_02520_),
    .A2(_02521_),
    .A3(_02524_),
    .A4(_02526_),
    .ZN(_02527_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08236_ (.A1(_02517_),
    .A2(_02527_),
    .ZN(_02528_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08237_ (.A1(_00749_),
    .A2(_00561_),
    .ZN(_02529_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _08238_ (.A1(_00936_),
    .A2(_00980_),
    .A3(_00964_),
    .ZN(_02530_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08239_ (.A1(_00798_),
    .A2(_02522_),
    .ZN(_02531_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _08240_ (.A1(_00836_),
    .A2(_02529_),
    .A3(_02530_),
    .A4(_02531_),
    .ZN(_02532_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _08241_ (.A1(_00934_),
    .A2(_00965_),
    .A3(_02525_),
    .ZN(_02533_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08242_ (.A1(_02532_),
    .A2(_02533_),
    .ZN(_02534_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _08243_ (.A1(_00780_),
    .A2(_00655_),
    .A3(_00574_),
    .ZN(_02535_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08244_ (.I(_02535_),
    .Z(_02536_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08245_ (.I(_02536_),
    .Z(_02537_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _08246_ (.A1(_00966_),
    .A2(_00681_),
    .A3(_02509_),
    .ZN(_02538_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08247_ (.A1(_00523_),
    .A2(_02537_),
    .B(_02538_),
    .ZN(_02539_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08248_ (.A1(_00912_),
    .A2(_00533_),
    .A3(_00981_),
    .A4(_01787_),
    .Z(_02540_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _08249_ (.A1(_00565_),
    .A2(_01927_),
    .A3(_02525_),
    .ZN(_02541_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08250_ (.A1(_01108_),
    .A2(_05746_),
    .ZN(_02542_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08251_ (.A1(_00726_),
    .A2(_02518_),
    .A3(_02542_),
    .ZN(_02543_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08252_ (.A1(_02537_),
    .A2(_02540_),
    .B(_02541_),
    .C(_02543_),
    .ZN(_02544_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08253_ (.A1(_02534_),
    .A2(_02539_),
    .A3(_02544_),
    .ZN(_02545_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08254_ (.A1(_02512_),
    .A2(_02528_),
    .A3(_02545_),
    .ZN(_02546_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08255_ (.I(_00968_),
    .Z(_02547_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08256_ (.I(_02547_),
    .Z(_02548_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08257_ (.I(_00535_),
    .Z(_02549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08258_ (.A1(_02146_),
    .A2(_02549_),
    .ZN(_02550_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08259_ (.I(net1),
    .Z(_02551_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08260_ (.I(_02551_),
    .Z(_02552_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08261_ (.I(_02552_),
    .Z(_02553_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08262_ (.I(_02553_),
    .Z(_02554_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08263_ (.I(_02554_),
    .Z(_02555_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08264_ (.A1(_05725_),
    .A2(_02339_),
    .Z(_02556_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08265_ (.I(_02556_),
    .Z(_02557_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08266_ (.A1(_02554_),
    .A2(_02557_),
    .ZN(_02558_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08267_ (.I(_01802_),
    .Z(_02559_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08268_ (.I(_02559_),
    .Z(_02560_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08269_ (.I(_02560_),
    .Z(_02561_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08270_ (.I(_02561_),
    .Z(_02562_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08271_ (.A1(_02484_),
    .A2(_02555_),
    .B(_02558_),
    .C(_02562_),
    .ZN(_02563_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08272_ (.I(_00563_),
    .Z(_02564_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08273_ (.I(_02564_),
    .Z(_02565_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08274_ (.I(_02565_),
    .Z(_02566_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08275_ (.I(_02566_),
    .Z(_02567_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08276_ (.A1(_02550_),
    .A2(_02563_),
    .B(_02567_),
    .ZN(_02568_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08277_ (.A1(_02548_),
    .A2(_02568_),
    .B(_02546_),
    .ZN(_02569_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08278_ (.I(_00882_),
    .Z(_02570_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08279_ (.A1(_02485_),
    .A2(_02546_),
    .B(_02569_),
    .C(_02570_),
    .ZN(_00119_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08280_ (.I(_02186_),
    .Z(_02571_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _08281_ (.A1(_02312_),
    .A2(_02175_),
    .A3(_02466_),
    .ZN(_02572_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08282_ (.I(_02572_),
    .Z(_02573_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08283_ (.I(_02573_),
    .Z(_02574_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08284_ (.I(_02572_),
    .Z(_02575_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08285_ (.A1(\as2650.stack[6][8] ),
    .A2(_02575_),
    .ZN(_02576_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08286_ (.A1(_02451_),
    .A2(_02191_),
    .A3(_02453_),
    .ZN(_02577_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08287_ (.I(_02577_),
    .Z(_02578_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08288_ (.I(_02578_),
    .Z(_02579_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08289_ (.A1(_02571_),
    .A2(_02574_),
    .B(_02576_),
    .C(_02579_),
    .ZN(_00120_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08290_ (.I(_02198_),
    .Z(_02580_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08291_ (.I(_02572_),
    .Z(_02581_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08292_ (.A1(\as2650.stack[6][9] ),
    .A2(_02581_),
    .ZN(_02582_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08293_ (.A1(_02580_),
    .A2(_02574_),
    .B(_02582_),
    .C(_02579_),
    .ZN(_00121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08294_ (.I(_02205_),
    .Z(_02583_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08295_ (.A1(\as2650.stack[6][10] ),
    .A2(_02581_),
    .ZN(_02584_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08296_ (.A1(_02583_),
    .A2(_02574_),
    .B(_02584_),
    .C(_02579_),
    .ZN(_00122_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08297_ (.I(_02211_),
    .Z(_02585_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08298_ (.A1(\as2650.stack[6][11] ),
    .A2(_02581_),
    .ZN(_02586_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08299_ (.A1(_02585_),
    .A2(_02574_),
    .B(_02586_),
    .C(_02579_),
    .ZN(_00123_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08300_ (.I(_02218_),
    .Z(_02587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08301_ (.I(_02573_),
    .Z(_02588_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08302_ (.A1(\as2650.stack[6][12] ),
    .A2(_02581_),
    .ZN(_02589_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08303_ (.I(_02578_),
    .Z(_02590_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08304_ (.A1(_02587_),
    .A2(_02588_),
    .B(_02589_),
    .C(_02590_),
    .ZN(_00124_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08305_ (.I(_02225_),
    .Z(_02591_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08306_ (.A1(\as2650.stack[6][13] ),
    .A2(_02573_),
    .ZN(_02592_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08307_ (.A1(_02591_),
    .A2(_02588_),
    .B(_02592_),
    .C(_02590_),
    .ZN(_00125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08308_ (.I(_02232_),
    .Z(_02593_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08309_ (.A1(\as2650.stack[6][14] ),
    .A2(_02573_),
    .ZN(_02594_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08310_ (.A1(_02593_),
    .A2(_02588_),
    .B(_02594_),
    .C(_02590_),
    .ZN(_00126_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _08311_ (.A1(_02312_),
    .A2(_01825_),
    .A3(_02466_),
    .ZN(_02595_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08312_ (.I(_02595_),
    .Z(_02596_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08313_ (.I(_02596_),
    .Z(_02597_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08314_ (.I(_02595_),
    .Z(_02598_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08315_ (.A1(\as2650.stack[5][8] ),
    .A2(_02598_),
    .ZN(_02599_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08316_ (.A1(_02451_),
    .A2(_01771_),
    .A3(_02453_),
    .ZN(_02600_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08317_ (.I(_02600_),
    .Z(_02601_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08318_ (.I(_02601_),
    .Z(_02602_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08319_ (.A1(_02571_),
    .A2(_02597_),
    .B(_02599_),
    .C(_02602_),
    .ZN(_00127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08320_ (.I(_02595_),
    .Z(_02603_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08321_ (.A1(\as2650.stack[5][9] ),
    .A2(_02603_),
    .ZN(_02604_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08322_ (.A1(_02580_),
    .A2(_02597_),
    .B(_02604_),
    .C(_02602_),
    .ZN(_00128_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08323_ (.A1(\as2650.stack[5][10] ),
    .A2(_02603_),
    .ZN(_02605_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08324_ (.A1(_02583_),
    .A2(_02597_),
    .B(_02605_),
    .C(_02602_),
    .ZN(_00129_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08325_ (.A1(\as2650.stack[5][11] ),
    .A2(_02603_),
    .ZN(_02606_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08326_ (.A1(_02585_),
    .A2(_02597_),
    .B(_02606_),
    .C(_02602_),
    .ZN(_00130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08327_ (.I(_02596_),
    .Z(_02607_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08328_ (.A1(\as2650.stack[5][12] ),
    .A2(_02603_),
    .ZN(_02608_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08329_ (.I(_02601_),
    .Z(_02609_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08330_ (.A1(_02587_),
    .A2(_02607_),
    .B(_02608_),
    .C(_02609_),
    .ZN(_00131_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08331_ (.A1(\as2650.stack[5][13] ),
    .A2(_02596_),
    .ZN(_02610_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08332_ (.A1(_02591_),
    .A2(_02607_),
    .B(_02610_),
    .C(_02609_),
    .ZN(_00132_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08333_ (.A1(\as2650.stack[5][14] ),
    .A2(_02596_),
    .ZN(_02611_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08334_ (.A1(_02593_),
    .A2(_02607_),
    .B(_02611_),
    .C(_02609_),
    .ZN(_00133_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _08335_ (.A1(_01772_),
    .A2(_02260_),
    .A3(_02466_),
    .ZN(_02612_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08336_ (.I(_02612_),
    .Z(_02613_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08337_ (.I(_02613_),
    .Z(_02614_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08338_ (.I(_02612_),
    .Z(_02615_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08339_ (.A1(\as2650.stack[4][8] ),
    .A2(_02615_),
    .ZN(_02616_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _08340_ (.A1(_02394_),
    .A2(_02401_),
    .ZN(_02617_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08341_ (.A1(_01767_),
    .A2(_02617_),
    .ZN(_02618_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08342_ (.I(_02618_),
    .Z(_02619_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08343_ (.I(_02619_),
    .Z(_02620_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08344_ (.A1(_02571_),
    .A2(_02614_),
    .B(_02616_),
    .C(_02620_),
    .ZN(_00134_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08345_ (.I(_02612_),
    .Z(_02621_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08346_ (.A1(\as2650.stack[4][9] ),
    .A2(_02621_),
    .ZN(_02622_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08347_ (.A1(_02580_),
    .A2(_02614_),
    .B(_02622_),
    .C(_02620_),
    .ZN(_00135_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08348_ (.A1(\as2650.stack[4][10] ),
    .A2(_02621_),
    .ZN(_02623_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08349_ (.A1(_02583_),
    .A2(_02614_),
    .B(_02623_),
    .C(_02620_),
    .ZN(_00136_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08350_ (.A1(\as2650.stack[4][11] ),
    .A2(_02621_),
    .ZN(_02624_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08351_ (.A1(_02585_),
    .A2(_02614_),
    .B(_02624_),
    .C(_02620_),
    .ZN(_00137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08352_ (.I(_02613_),
    .Z(_02625_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08353_ (.A1(\as2650.stack[4][12] ),
    .A2(_02621_),
    .ZN(_02626_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08354_ (.I(_02619_),
    .Z(_02627_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08355_ (.A1(_02587_),
    .A2(_02625_),
    .B(_02626_),
    .C(_02627_),
    .ZN(_00138_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08356_ (.A1(\as2650.stack[4][13] ),
    .A2(_02613_),
    .ZN(_02628_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08357_ (.A1(_02591_),
    .A2(_02625_),
    .B(_02628_),
    .C(_02627_),
    .ZN(_00139_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08358_ (.A1(\as2650.stack[4][14] ),
    .A2(_02613_),
    .ZN(_02629_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08359_ (.A1(_02593_),
    .A2(_02625_),
    .B(_02629_),
    .C(_02627_),
    .ZN(_00140_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08360_ (.I(_01761_),
    .Z(_02630_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08361_ (.I(_02300_),
    .Z(_02631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08362_ (.I(_02631_),
    .Z(_02632_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _08363_ (.A1(_01783_),
    .A2(_01785_),
    .A3(_02399_),
    .A4(_01807_),
    .ZN(_02633_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08364_ (.I(_02633_),
    .Z(_02634_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08365_ (.A1(\as2650.stack[12][0] ),
    .A2(_02634_),
    .ZN(_02635_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08366_ (.A1(_02259_),
    .A2(_02307_),
    .B(_02309_),
    .ZN(_02636_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08367_ (.A1(_02630_),
    .A2(_02632_),
    .B1(_02635_),
    .B2(_02636_),
    .ZN(_00141_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08368_ (.I(_01846_),
    .Z(_02637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08369_ (.A1(\as2650.stack[12][1] ),
    .A2(_02634_),
    .ZN(_02638_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08370_ (.I(_02293_),
    .Z(_02639_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08371_ (.I(_02301_),
    .Z(_02640_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08372_ (.A1(_02268_),
    .A2(_02639_),
    .B(_02640_),
    .ZN(_02641_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08373_ (.A1(_02637_),
    .A2(_02632_),
    .B1(_02638_),
    .B2(_02641_),
    .ZN(_00142_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08374_ (.I(_01862_),
    .Z(_02642_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08375_ (.A1(\as2650.stack[12][2] ),
    .A2(_02634_),
    .ZN(_02643_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08376_ (.A1(_02273_),
    .A2(_02639_),
    .B(_02640_),
    .ZN(_02644_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08377_ (.A1(_02642_),
    .A2(_02632_),
    .B1(_02643_),
    .B2(_02644_),
    .ZN(_00143_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08378_ (.I(_01873_),
    .Z(_02645_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08379_ (.A1(\as2650.stack[12][3] ),
    .A2(_02634_),
    .ZN(_02646_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08380_ (.A1(_02276_),
    .A2(_02639_),
    .B(_02640_),
    .ZN(_02647_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08381_ (.A1(_02645_),
    .A2(_02632_),
    .B1(_02646_),
    .B2(_02647_),
    .ZN(_00144_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08382_ (.I(_01883_),
    .Z(_02648_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08383_ (.I(_02301_),
    .Z(_02649_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08384_ (.I(_02633_),
    .Z(_02650_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08385_ (.A1(\as2650.stack[12][4] ),
    .A2(_02650_),
    .ZN(_02651_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08386_ (.A1(_02281_),
    .A2(_02639_),
    .B(_02640_),
    .ZN(_02652_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08387_ (.A1(_02648_),
    .A2(_02649_),
    .B1(_02651_),
    .B2(_02652_),
    .ZN(_00145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08388_ (.I(_01895_),
    .Z(_02653_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08389_ (.A1(\as2650.stack[12][5] ),
    .A2(_02650_),
    .ZN(_02654_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08390_ (.A1(_02284_),
    .A2(_02296_),
    .B(_02631_),
    .ZN(_02655_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08391_ (.A1(_02653_),
    .A2(_02649_),
    .B1(_02654_),
    .B2(_02655_),
    .ZN(_00146_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08392_ (.I(_01908_),
    .Z(_02656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08393_ (.A1(\as2650.stack[12][6] ),
    .A2(_02650_),
    .ZN(_02657_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08394_ (.A1(_02288_),
    .A2(_02296_),
    .B(_02631_),
    .ZN(_02658_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08395_ (.A1(_02656_),
    .A2(_02649_),
    .B1(_02657_),
    .B2(_02658_),
    .ZN(_00147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08396_ (.I(_01918_),
    .Z(_02659_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08397_ (.A1(\as2650.stack[12][7] ),
    .A2(_02650_),
    .ZN(_02660_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08398_ (.A1(_02291_),
    .A2(_02296_),
    .B(_02631_),
    .ZN(_02661_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08399_ (.A1(_02659_),
    .A2(_02649_),
    .B1(_02660_),
    .B2(_02661_),
    .ZN(_00148_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08400_ (.A1(_02444_),
    .A2(_02617_),
    .ZN(_02662_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08401_ (.I(_02662_),
    .Z(_02663_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08402_ (.I(_02663_),
    .Z(_02664_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08403_ (.I(_02662_),
    .Z(_02665_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08404_ (.A1(\as2650.stack[3][8] ),
    .A2(_02665_),
    .ZN(_02666_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08405_ (.I(_01766_),
    .Z(_02667_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08406_ (.A1(_02667_),
    .A2(_02318_),
    .A3(_02408_),
    .ZN(_02668_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08407_ (.I(_02668_),
    .Z(_02669_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08408_ (.I(_02669_),
    .Z(_02670_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08409_ (.A1(_02571_),
    .A2(_02664_),
    .B(_02666_),
    .C(_02670_),
    .ZN(_00149_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08410_ (.I(_02662_),
    .Z(_02671_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08411_ (.A1(\as2650.stack[3][9] ),
    .A2(_02671_),
    .ZN(_02672_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08412_ (.A1(_02580_),
    .A2(_02664_),
    .B(_02672_),
    .C(_02670_),
    .ZN(_00150_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08413_ (.A1(\as2650.stack[3][10] ),
    .A2(_02671_),
    .ZN(_02673_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08414_ (.A1(_02583_),
    .A2(_02664_),
    .B(_02673_),
    .C(_02670_),
    .ZN(_00151_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08415_ (.A1(\as2650.stack[3][11] ),
    .A2(_02671_),
    .ZN(_02674_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08416_ (.A1(_02585_),
    .A2(_02664_),
    .B(_02674_),
    .C(_02670_),
    .ZN(_00152_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08417_ (.I(_02663_),
    .Z(_02675_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08418_ (.A1(\as2650.stack[3][12] ),
    .A2(_02671_),
    .ZN(_02676_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08419_ (.I(_02669_),
    .Z(_02677_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08420_ (.A1(_02587_),
    .A2(_02675_),
    .B(_02676_),
    .C(_02677_),
    .ZN(_00153_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08421_ (.A1(\as2650.stack[3][13] ),
    .A2(_02663_),
    .ZN(_02678_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08422_ (.A1(_02591_),
    .A2(_02675_),
    .B(_02678_),
    .C(_02677_),
    .ZN(_00154_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08423_ (.A1(\as2650.stack[3][14] ),
    .A2(_02663_),
    .ZN(_02679_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08424_ (.A1(_02593_),
    .A2(_02675_),
    .B(_02679_),
    .C(_02677_),
    .ZN(_00155_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08425_ (.I(_02186_),
    .Z(_02680_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _08426_ (.A1(_01821_),
    .A2(_02175_),
    .A3(_02408_),
    .ZN(_02681_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08427_ (.I(_02681_),
    .Z(_02682_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08428_ (.I(_02682_),
    .Z(_02683_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08429_ (.I(_02681_),
    .Z(_02684_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08430_ (.A1(\as2650.stack[2][8] ),
    .A2(_02684_),
    .ZN(_02685_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08431_ (.A1(_02667_),
    .A2(_02191_),
    .A3(_02407_),
    .ZN(_02686_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08432_ (.I(_02686_),
    .Z(_02687_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08433_ (.I(_02687_),
    .Z(_02688_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08434_ (.A1(_02680_),
    .A2(_02683_),
    .B(_02685_),
    .C(_02688_),
    .ZN(_00156_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08435_ (.I(_02198_),
    .Z(_02689_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08436_ (.I(_02681_),
    .Z(_02690_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08437_ (.A1(\as2650.stack[2][9] ),
    .A2(_02690_),
    .ZN(_02691_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08438_ (.A1(_02689_),
    .A2(_02683_),
    .B(_02691_),
    .C(_02688_),
    .ZN(_00157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08439_ (.I(_02205_),
    .Z(_02692_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08440_ (.A1(\as2650.stack[2][10] ),
    .A2(_02690_),
    .ZN(_02693_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08441_ (.A1(_02692_),
    .A2(_02683_),
    .B(_02693_),
    .C(_02688_),
    .ZN(_00158_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08442_ (.I(_02211_),
    .Z(_02694_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08443_ (.A1(\as2650.stack[2][11] ),
    .A2(_02690_),
    .ZN(_02695_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08444_ (.A1(_02694_),
    .A2(_02683_),
    .B(_02695_),
    .C(_02688_),
    .ZN(_00159_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08445_ (.I(_02218_),
    .Z(_02696_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08446_ (.I(_02682_),
    .Z(_02697_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08447_ (.A1(\as2650.stack[2][12] ),
    .A2(_02690_),
    .ZN(_02698_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08448_ (.I(_02687_),
    .Z(_02699_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08449_ (.A1(_02696_),
    .A2(_02697_),
    .B(_02698_),
    .C(_02699_),
    .ZN(_00160_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08450_ (.I(_02225_),
    .Z(_02700_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08451_ (.A1(\as2650.stack[2][13] ),
    .A2(_02682_),
    .ZN(_02701_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08452_ (.A1(_02700_),
    .A2(_02697_),
    .B(_02701_),
    .C(_02699_),
    .ZN(_00161_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08453_ (.I(_02232_),
    .Z(_02702_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08454_ (.A1(\as2650.stack[2][14] ),
    .A2(_02682_),
    .ZN(_02703_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08455_ (.A1(_02702_),
    .A2(_02697_),
    .B(_02703_),
    .C(_02699_),
    .ZN(_00162_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _08456_ (.A1(_01821_),
    .A2(_01825_),
    .A3(_02408_),
    .ZN(_02704_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08457_ (.I(_02704_),
    .Z(_02705_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08458_ (.I(_02705_),
    .Z(_02706_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08459_ (.I(_02704_),
    .Z(_02707_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08460_ (.A1(\as2650.stack[1][8] ),
    .A2(_02707_),
    .ZN(_02708_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08461_ (.A1(_02667_),
    .A2(_01771_),
    .A3(_02407_),
    .ZN(_02709_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08462_ (.I(_02709_),
    .Z(_02710_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08463_ (.I(_02710_),
    .Z(_02711_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08464_ (.A1(_02680_),
    .A2(_02706_),
    .B(_02708_),
    .C(_02711_),
    .ZN(_00163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08465_ (.I(_02704_),
    .Z(_02712_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08466_ (.A1(\as2650.stack[1][9] ),
    .A2(_02712_),
    .ZN(_02713_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08467_ (.A1(_02689_),
    .A2(_02706_),
    .B(_02713_),
    .C(_02711_),
    .ZN(_00164_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08468_ (.A1(\as2650.stack[1][10] ),
    .A2(_02712_),
    .ZN(_02714_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08469_ (.A1(_02692_),
    .A2(_02706_),
    .B(_02714_),
    .C(_02711_),
    .ZN(_00165_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08470_ (.A1(\as2650.stack[1][11] ),
    .A2(_02712_),
    .ZN(_02715_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08471_ (.A1(_02694_),
    .A2(_02706_),
    .B(_02715_),
    .C(_02711_),
    .ZN(_00166_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08472_ (.I(_02705_),
    .Z(_02716_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08473_ (.A1(\as2650.stack[1][12] ),
    .A2(_02712_),
    .ZN(_02717_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08474_ (.I(_02710_),
    .Z(_02718_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08475_ (.A1(_02696_),
    .A2(_02716_),
    .B(_02717_),
    .C(_02718_),
    .ZN(_00167_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08476_ (.A1(\as2650.stack[1][13] ),
    .A2(_02705_),
    .ZN(_02719_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08477_ (.A1(_02700_),
    .A2(_02716_),
    .B(_02719_),
    .C(_02718_),
    .ZN(_00168_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08478_ (.A1(\as2650.stack[1][14] ),
    .A2(_02705_),
    .ZN(_02720_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08479_ (.A1(_02702_),
    .A2(_02716_),
    .B(_02720_),
    .C(_02718_),
    .ZN(_00169_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08480_ (.A1(_02444_),
    .A2(_02395_),
    .ZN(_02721_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08481_ (.I(_02721_),
    .Z(_02722_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08482_ (.I(_02722_),
    .Z(_02723_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08483_ (.I(_02721_),
    .Z(_02724_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08484_ (.A1(\as2650.stack[15][8] ),
    .A2(_02724_),
    .ZN(_02725_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08485_ (.A1(_02667_),
    .A2(_01778_),
    .A3(_02318_),
    .ZN(_02726_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08486_ (.I(_02726_),
    .Z(_02727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08487_ (.I(_02727_),
    .Z(_02728_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08488_ (.A1(_02680_),
    .A2(_02723_),
    .B(_02725_),
    .C(_02728_),
    .ZN(_00170_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08489_ (.I(_02721_),
    .Z(_02729_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08490_ (.A1(\as2650.stack[15][9] ),
    .A2(_02729_),
    .ZN(_02730_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08491_ (.A1(_02689_),
    .A2(_02723_),
    .B(_02730_),
    .C(_02728_),
    .ZN(_00171_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08492_ (.A1(\as2650.stack[15][10] ),
    .A2(_02729_),
    .ZN(_02731_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08493_ (.A1(_02692_),
    .A2(_02723_),
    .B(_02731_),
    .C(_02728_),
    .ZN(_00172_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08494_ (.A1(\as2650.stack[15][11] ),
    .A2(_02729_),
    .ZN(_02732_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08495_ (.A1(_02694_),
    .A2(_02723_),
    .B(_02732_),
    .C(_02728_),
    .ZN(_00173_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08496_ (.I(_02722_),
    .Z(_02733_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08497_ (.A1(\as2650.stack[15][12] ),
    .A2(_02729_),
    .ZN(_02734_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08498_ (.I(_02727_),
    .Z(_02735_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08499_ (.A1(_02696_),
    .A2(_02733_),
    .B(_02734_),
    .C(_02735_),
    .ZN(_00174_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08500_ (.A1(\as2650.stack[15][13] ),
    .A2(_02722_),
    .ZN(_02736_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08501_ (.A1(_02700_),
    .A2(_02733_),
    .B(_02736_),
    .C(_02735_),
    .ZN(_00175_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08502_ (.A1(\as2650.stack[15][14] ),
    .A2(_02722_),
    .ZN(_02737_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08503_ (.A1(_02702_),
    .A2(_02733_),
    .B(_02737_),
    .C(_02735_),
    .ZN(_00176_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08504_ (.I(_00672_),
    .Z(_02738_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08505_ (.I(_01802_),
    .Z(_02739_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _08506_ (.A1(_02738_),
    .A2(_02739_),
    .ZN(_02740_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08507_ (.I(_00940_),
    .Z(_02741_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08508_ (.A1(_00582_),
    .A2(_02741_),
    .B1(_02334_),
    .B2(_02556_),
    .ZN(_02742_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08509_ (.I(_02742_),
    .ZN(_02743_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08510_ (.I(_02507_),
    .Z(_02744_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _08511_ (.A1(_00944_),
    .A2(_02740_),
    .B1(_02743_),
    .B2(_02744_),
    .ZN(_02745_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _08512_ (.A1(_00782_),
    .A2(_00894_),
    .A3(_00967_),
    .A4(_00544_),
    .ZN(_02746_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08513_ (.I(_02564_),
    .Z(_02747_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08514_ (.I(_01018_),
    .Z(_02748_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08515_ (.I(_00982_),
    .Z(_02749_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08516_ (.I(_02739_),
    .Z(_02750_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _08517_ (.A1(_02747_),
    .A2(_00571_),
    .A3(_02748_),
    .B1(_02749_),
    .B2(_02750_),
    .ZN(_02751_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08518_ (.A1(_02744_),
    .A2(_02751_),
    .ZN(_02752_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08519_ (.A1(_02745_),
    .A2(_02746_),
    .A3(_02752_),
    .ZN(_02753_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _08520_ (.A1(_00913_),
    .A2(_00918_),
    .A3(_02749_),
    .A4(_01787_),
    .ZN(_02754_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08521_ (.A1(_00625_),
    .A2(_00824_),
    .B(_00904_),
    .ZN(_02755_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08522_ (.A1(_02740_),
    .A2(_02755_),
    .ZN(_02756_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08523_ (.A1(_02738_),
    .A2(_01764_),
    .ZN(_02757_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _08524_ (.A1(_00972_),
    .A2(_00813_),
    .A3(_00955_),
    .B(_02738_),
    .ZN(_02758_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08525_ (.A1(_00502_),
    .A2(_02492_),
    .B(_02757_),
    .C(_02758_),
    .ZN(_02759_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08526_ (.A1(_00918_),
    .A2(_00979_),
    .B(_02759_),
    .ZN(_02760_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08527_ (.I(_01793_),
    .Z(_02761_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08528_ (.I(_00551_),
    .Z(_02762_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _08529_ (.A1(_00581_),
    .A2(_02564_),
    .A3(_00671_),
    .ZN(_02763_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _08530_ (.A1(_00959_),
    .A2(_02747_),
    .B1(_02761_),
    .B2(_02762_),
    .C(_02763_),
    .ZN(_02764_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _08531_ (.A1(_02754_),
    .A2(_02756_),
    .A3(_02760_),
    .A4(_02764_),
    .ZN(_02765_));
 gf180mcu_fd_sc_mcu7t5v0__oai33_1 _08532_ (.A1(_00791_),
    .A2(_02564_),
    .A3(_01063_),
    .B1(_02761_),
    .B2(_02492_),
    .B3(_00896_),
    .ZN(_02766_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08533_ (.A1(_00581_),
    .A2(_00949_),
    .ZN(_02767_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08534_ (.I(_02767_),
    .ZN(_02768_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _08535_ (.A1(_02762_),
    .A2(_00955_),
    .A3(_00822_),
    .A4(_02768_),
    .ZN(_02769_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _08536_ (.A1(_00913_),
    .A2(_02347_),
    .A3(_02761_),
    .A4(_02339_),
    .ZN(_02770_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08537_ (.A1(_00804_),
    .A2(_00552_),
    .A3(_02516_),
    .ZN(_02771_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08538_ (.A1(_00815_),
    .A2(_02769_),
    .B(_02770_),
    .C(_02771_),
    .ZN(_02772_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08539_ (.A1(_02766_),
    .A2(_02772_),
    .ZN(_02773_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08540_ (.A1(_00912_),
    .A2(_02491_),
    .A3(_02513_),
    .A4(_00700_),
    .Z(_02774_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _08541_ (.A1(_01108_),
    .A2(_00826_),
    .A3(_02498_),
    .A4(_02774_),
    .ZN(_02775_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08542_ (.A1(_00534_),
    .A2(_00813_),
    .A3(_00564_),
    .ZN(_02776_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08543_ (.A1(_02773_),
    .A2(_02775_),
    .A3(_02776_),
    .ZN(_02777_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _08544_ (.A1(_02753_),
    .A2(_02765_),
    .A3(_02777_),
    .ZN(_02778_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08545_ (.A1(_01271_),
    .A2(_01208_),
    .A3(_01053_),
    .ZN(_02779_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _08546_ (.A1(_01615_),
    .A2(_01533_),
    .A3(_01420_),
    .A4(_01324_),
    .ZN(_02780_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08547_ (.A1(_02779_),
    .A2(_02780_),
    .ZN(_02781_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08548_ (.I(_01703_),
    .Z(_02782_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08549_ (.A1(_02782_),
    .A2(_00817_),
    .ZN(_02783_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08550_ (.I(_01618_),
    .Z(_02784_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08551_ (.A1(_02784_),
    .A2(_00956_),
    .A3(_01697_),
    .ZN(_02785_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08552_ (.A1(_02781_),
    .A2(_02783_),
    .B(_02785_),
    .ZN(_02786_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08553_ (.A1(_01139_),
    .A2(_01188_),
    .A3(_01304_),
    .A4(_01373_),
    .Z(_02787_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08554_ (.A1(_01461_),
    .A2(_02787_),
    .ZN(_02788_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08555_ (.A1(_01013_),
    .A2(_01694_),
    .ZN(_02789_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _08556_ (.A1(_01514_),
    .A2(_01606_),
    .A3(_02788_),
    .B(_02789_),
    .ZN(_02790_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08557_ (.A1(_01442_),
    .A2(_01443_),
    .Z(_02791_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08558_ (.A1(_01679_),
    .A2(_01689_),
    .ZN(_02792_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08559_ (.A1(_01594_),
    .A2(_02792_),
    .ZN(_02793_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08560_ (.A1(_02791_),
    .A2(_01498_),
    .A3(_02793_),
    .ZN(_02794_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08561_ (.A1(_01125_),
    .A2(_01176_),
    .A3(_01287_),
    .A4(_01358_),
    .Z(_02795_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08562_ (.A1(_01676_),
    .A2(_01677_),
    .ZN(_02796_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08563_ (.A1(_01672_),
    .A2(_02796_),
    .ZN(_02797_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _08564_ (.A1(_01350_),
    .A2(_01180_),
    .A3(_01601_),
    .ZN(_02798_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08565_ (.A1(_01450_),
    .A2(_01356_),
    .ZN(_02799_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08566_ (.A1(_01169_),
    .A2(_01170_),
    .B(_01176_),
    .ZN(_02800_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08567_ (.A1(_01289_),
    .A2(_02800_),
    .B(_01294_),
    .ZN(_02801_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08568_ (.A1(_01364_),
    .A2(_02801_),
    .B(_01358_),
    .ZN(_02802_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _08569_ (.A1(_02799_),
    .A2(_02802_),
    .Z(_02803_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08570_ (.I(_02803_),
    .ZN(_02804_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08571_ (.A1(_01498_),
    .A2(_01500_),
    .ZN(_02805_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08572_ (.A1(_01595_),
    .A2(_02805_),
    .B(_01594_),
    .ZN(_02806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08573_ (.A1(_01682_),
    .A2(_02806_),
    .ZN(_02807_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08574_ (.A1(_02792_),
    .A2(_02807_),
    .ZN(_02808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08575_ (.A1(_02797_),
    .A2(_02808_),
    .ZN(_02809_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08576_ (.A1(_01845_),
    .A2(_01681_),
    .B1(_02804_),
    .B2(_02794_),
    .C(_02809_),
    .ZN(_02810_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08577_ (.A1(_02798_),
    .A2(_02810_),
    .ZN(_02811_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _08578_ (.A1(net79),
    .A2(_02792_),
    .A3(_02797_),
    .B(_02811_),
    .ZN(_02812_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08579_ (.A1(_02794_),
    .A2(_02795_),
    .B(_02812_),
    .ZN(_02813_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08580_ (.A1(_00795_),
    .A2(_02813_),
    .ZN(_02814_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08581_ (.A1(_00538_),
    .A2(_02786_),
    .B1(_02790_),
    .B2(_02814_),
    .ZN(_02815_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08582_ (.I(_00839_),
    .Z(_02816_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08583_ (.I(_01942_),
    .Z(_02817_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08584_ (.I(_02817_),
    .Z(_02818_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08585_ (.I(_01947_),
    .Z(_02819_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08586_ (.I(_01810_),
    .Z(_02820_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08587_ (.I(_01953_),
    .Z(_02821_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08588_ (.A1(\as2650.stack[8][6] ),
    .A2(_02820_),
    .B1(_02821_),
    .B2(\as2650.stack[9][6] ),
    .ZN(_02822_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08589_ (.I(_01939_),
    .Z(_02823_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08590_ (.I(_02823_),
    .Z(_02824_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08591_ (.A1(\as2650.stack[11][6] ),
    .A2(_02824_),
    .B1(_01964_),
    .B2(\as2650.stack[10][6] ),
    .ZN(_02825_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08592_ (.A1(_02819_),
    .A2(_02822_),
    .A3(_02825_),
    .ZN(_02826_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08593_ (.I(_01946_),
    .Z(_02827_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08594_ (.I(_02823_),
    .Z(_02828_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08595_ (.I(_01963_),
    .Z(_02829_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08596_ (.A1(\as2650.stack[15][6] ),
    .A2(_02828_),
    .B1(_02829_),
    .B2(\as2650.stack[14][6] ),
    .ZN(_02830_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08597_ (.A1(\as2650.stack[12][6] ),
    .A2(_02820_),
    .B1(_02821_),
    .B2(\as2650.stack[13][6] ),
    .ZN(_02831_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08598_ (.A1(_02827_),
    .A2(_02830_),
    .A3(_02831_),
    .ZN(_02832_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08599_ (.A1(_02826_),
    .A2(_02832_),
    .ZN(_02833_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08600_ (.I(_01947_),
    .Z(_02834_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08601_ (.I(_01810_),
    .Z(_02835_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08602_ (.A1(\as2650.stack[0][6] ),
    .A2(_02835_),
    .B1(_01954_),
    .B2(\as2650.stack[1][6] ),
    .ZN(_02836_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08603_ (.I(_01940_),
    .Z(_02837_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08604_ (.I(_01963_),
    .Z(_02838_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08605_ (.A1(\as2650.stack[3][6] ),
    .A2(_02837_),
    .B1(_02838_),
    .B2(\as2650.stack[2][6] ),
    .ZN(_02839_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08606_ (.A1(_02834_),
    .A2(_02836_),
    .A3(_02839_),
    .ZN(_02840_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08607_ (.A1(\as2650.stack[7][6] ),
    .A2(_02837_),
    .B1(_02838_),
    .B2(\as2650.stack[6][6] ),
    .ZN(_02841_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08608_ (.I(_01953_),
    .Z(_02842_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08609_ (.A1(\as2650.stack[4][6] ),
    .A2(_02835_),
    .B1(_02842_),
    .B2(\as2650.stack[5][6] ),
    .ZN(_02843_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08610_ (.A1(_02827_),
    .A2(_02841_),
    .A3(_02843_),
    .ZN(_02844_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08611_ (.A1(_02840_),
    .A2(_02844_),
    .B(_01943_),
    .ZN(_02845_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08612_ (.A1(_02818_),
    .A2(_02833_),
    .B(_02845_),
    .ZN(_02846_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _08613_ (.I(_02846_),
    .ZN(_02847_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08614_ (.I(_00897_),
    .Z(_02848_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08615_ (.I(_01426_),
    .Z(_02849_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08616_ (.I(_02849_),
    .Z(_02850_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08617_ (.I(_01623_),
    .Z(_02851_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08618_ (.I(_02851_),
    .Z(_02852_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08619_ (.I(_02852_),
    .Z(_02853_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08620_ (.I(_02853_),
    .Z(_02854_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08621_ (.A1(_02850_),
    .A2(_02554_),
    .A3(_02854_),
    .ZN(_02855_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08622_ (.I(_01080_),
    .Z(_02856_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08623_ (.I(_02856_),
    .Z(_02857_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08624_ (.I(_01216_),
    .Z(_02858_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08625_ (.I(_01265_),
    .Z(_02859_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08626_ (.I(_02859_),
    .Z(_02860_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08627_ (.I(net11),
    .Z(_02861_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08628_ (.I(_02861_),
    .Z(_02862_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08629_ (.I(_02862_),
    .Z(_02863_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08630_ (.I(_02863_),
    .Z(_02864_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08631_ (.I(_02864_),
    .Z(_02865_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _08632_ (.A1(_02857_),
    .A2(_02858_),
    .A3(_02860_),
    .A4(_02865_),
    .ZN(_02866_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08633_ (.A1(_02855_),
    .A2(_02866_),
    .B(_00851_),
    .ZN(_02867_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08634_ (.I(_00684_),
    .Z(_02868_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08635_ (.I(_02868_),
    .Z(_02869_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08636_ (.A1(_02869_),
    .A2(_01070_),
    .ZN(_02870_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08637_ (.A1(_01921_),
    .A2(_02781_),
    .B(_02488_),
    .ZN(_02871_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08638_ (.A1(_01911_),
    .A2(_02488_),
    .B(_02871_),
    .ZN(_02872_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08639_ (.A1(net101),
    .A2(_02852_),
    .B(_02494_),
    .C(_02750_),
    .ZN(_02873_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08640_ (.A1(_02853_),
    .A2(_02496_),
    .B(_02873_),
    .ZN(_02874_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08641_ (.A1(_05733_),
    .A2(_02337_),
    .ZN(_02875_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08642_ (.I(_01061_),
    .Z(_02876_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08643_ (.I(_02876_),
    .Z(_02877_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08644_ (.A1(_00536_),
    .A2(_02872_),
    .B1(_02874_),
    .B2(_02875_),
    .C(_02877_),
    .ZN(_02878_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08645_ (.I(_00962_),
    .Z(_02879_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08646_ (.A1(_01534_),
    .A2(_02876_),
    .ZN(_02880_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08647_ (.A1(_02879_),
    .A2(_02880_),
    .ZN(_02881_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _08648_ (.A1(_01609_),
    .A2(_02870_),
    .B(_02878_),
    .C(_02881_),
    .ZN(_02882_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08649_ (.I(_01704_),
    .Z(_02883_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08650_ (.I(_01581_),
    .Z(_02884_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08651_ (.I(_01499_),
    .Z(_02885_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08652_ (.A1(_02884_),
    .A2(_01617_),
    .A3(_02885_),
    .ZN(_02886_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08653_ (.A1(_02784_),
    .A2(_05851_),
    .A3(_02886_),
    .ZN(_02887_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08654_ (.I(_00897_),
    .Z(_02888_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _08655_ (.A1(_00963_),
    .A2(_02883_),
    .A3(_02887_),
    .B(_02888_),
    .ZN(_02889_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08656_ (.A1(_02848_),
    .A2(_02867_),
    .B1(_02882_),
    .B2(_02889_),
    .ZN(_02890_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08657_ (.I(_02490_),
    .Z(_02891_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08658_ (.A1(_02816_),
    .A2(_02847_),
    .B1(_02890_),
    .B2(_02891_),
    .ZN(_02892_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08659_ (.A1(_00807_),
    .A2(_02815_),
    .B(_02892_),
    .ZN(_02893_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08660_ (.A1(net53),
    .A2(_02778_),
    .B(_00883_),
    .ZN(_02894_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08661_ (.A1(_02778_),
    .A2(_02893_),
    .B(_02894_),
    .ZN(_00177_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08662_ (.A1(_05722_),
    .A2(_02778_),
    .B(_00846_),
    .ZN(_02895_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08663_ (.I(_01067_),
    .Z(_02896_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _08664_ (.A1(_02896_),
    .A2(_00817_),
    .B(_02783_),
    .C(_02562_),
    .ZN(_02897_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08665_ (.A1(_02562_),
    .A2(_02812_),
    .ZN(_02898_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08666_ (.A1(_02789_),
    .A2(_02898_),
    .ZN(_02899_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08667_ (.A1(_02897_),
    .A2(_02899_),
    .B(_00553_),
    .ZN(_02900_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08668_ (.I(_00529_),
    .Z(_02901_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08669_ (.I(_02901_),
    .Z(_02902_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08670_ (.I(_02902_),
    .Z(_02903_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08671_ (.I(_00670_),
    .Z(_02904_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08672_ (.I(_02904_),
    .Z(_02905_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08673_ (.A1(_00849_),
    .A2(_02505_),
    .ZN(_02906_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08674_ (.A1(_02862_),
    .A2(_01261_),
    .B1(_01072_),
    .B2(_01214_),
    .ZN(_02907_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08675_ (.I(_02907_),
    .ZN(_02908_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08676_ (.A1(_01624_),
    .A2(_01581_),
    .B1(_01211_),
    .B2(_01265_),
    .C(_02908_),
    .ZN(_02909_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08677_ (.I(_00600_),
    .Z(_02910_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08678_ (.A1(_00943_),
    .A2(_00500_),
    .A3(_02495_),
    .ZN(_02911_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _08679_ (.A1(_02910_),
    .A2(_01067_),
    .B1(_01522_),
    .B2(_02553_),
    .C(_02911_),
    .ZN(_02912_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08680_ (.A1(_01425_),
    .A2(_01499_),
    .B1(_01224_),
    .B2(_01080_),
    .ZN(_02913_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08681_ (.A1(_02909_),
    .A2(_02912_),
    .A3(_02913_),
    .Z(_02914_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _08682_ (.I(_01425_),
    .ZN(_02915_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08683_ (.A1(_01844_),
    .A2(_01215_),
    .B1(_01623_),
    .B2(_05735_),
    .ZN(_02916_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _08684_ (.A1(_01007_),
    .A2(_02915_),
    .B1(_01536_),
    .B2(net52),
    .C(_02916_),
    .ZN(_02917_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08685_ (.A1(_01760_),
    .A2(_01080_),
    .B1(_02862_),
    .B2(_01872_),
    .ZN(_02918_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08686_ (.A1(_05727_),
    .A2(_02910_),
    .B1(_01265_),
    .B2(_01861_),
    .ZN(_02919_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08687_ (.A1(_02911_),
    .A2(_02918_),
    .A3(_02919_),
    .ZN(_02920_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _08688_ (.A1(_01350_),
    .A2(_00625_),
    .A3(_00469_),
    .A4(_02338_),
    .ZN(_02921_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08689_ (.A1(_02917_),
    .A2(_02920_),
    .B(_02921_),
    .ZN(_02922_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _08690_ (.I(net29),
    .ZN(_02923_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _08691_ (.I(net10),
    .ZN(_02924_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08692_ (.I(_02924_),
    .Z(_02925_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08693_ (.A1(_01773_),
    .A2(_02925_),
    .B1(_02915_),
    .B2(net74),
    .ZN(_02926_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08694_ (.A1(_02173_),
    .A2(_01079_),
    .B1(_01215_),
    .B2(_01769_),
    .C(_02926_),
    .ZN(_02927_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _08695_ (.A1(_01776_),
    .A2(_01328_),
    .B1(_01536_),
    .B2(_02484_),
    .C(_02927_),
    .ZN(_02928_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _08696_ (.A1(_02923_),
    .A2(_02851_),
    .B1(_02346_),
    .B2(_00848_),
    .C(_02928_),
    .ZN(_02929_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08697_ (.A1(_02347_),
    .A2(_02494_),
    .A3(_02875_),
    .ZN(_02930_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _08698_ (.A1(_02914_),
    .A2(_02922_),
    .B1(_02929_),
    .B2(_02921_),
    .C(_02930_),
    .ZN(_02931_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _08699_ (.I(_02910_),
    .Z(_02932_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08700_ (.A1(_05722_),
    .A2(_02932_),
    .A3(_02930_),
    .ZN(_02933_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08701_ (.A1(_02497_),
    .A2(_02933_),
    .ZN(_02934_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08702_ (.A1(_05722_),
    .A2(_02906_),
    .B1(_02931_),
    .B2(_02934_),
    .ZN(_02935_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08703_ (.A1(_00793_),
    .A2(_02935_),
    .B(_02345_),
    .ZN(_02936_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08704_ (.A1(_02869_),
    .A2(_02936_),
    .ZN(_02937_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08705_ (.I(_02904_),
    .Z(_02938_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08706_ (.A1(_02880_),
    .A2(_02937_),
    .B(_02938_),
    .ZN(_02939_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08707_ (.A1(_02905_),
    .A2(_02883_),
    .B(_02939_),
    .ZN(_02940_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08708_ (.I(_00602_),
    .Z(_02941_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08709_ (.I(_02941_),
    .Z(_02942_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08710_ (.A1(_02942_),
    .A2(_02902_),
    .ZN(_02943_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08711_ (.A1(_02903_),
    .A2(_02940_),
    .B(_02943_),
    .ZN(_02944_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08712_ (.A1(_02891_),
    .A2(_02944_),
    .ZN(_02945_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08713_ (.I(_01942_),
    .Z(_02946_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08714_ (.A1(\as2650.stack[8][7] ),
    .A2(_01811_),
    .B1(_02842_),
    .B2(\as2650.stack[9][7] ),
    .ZN(_02947_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08715_ (.A1(\as2650.stack[11][7] ),
    .A2(_02837_),
    .B1(_02838_),
    .B2(\as2650.stack[10][7] ),
    .ZN(_02948_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08716_ (.A1(_02834_),
    .A2(_02947_),
    .A3(_02948_),
    .ZN(_02949_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08717_ (.I(_01946_),
    .Z(_02950_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08718_ (.I(_01940_),
    .Z(_02951_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08719_ (.A1(\as2650.stack[15][7] ),
    .A2(_02951_),
    .B1(_02838_),
    .B2(\as2650.stack[14][7] ),
    .ZN(_02952_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08720_ (.A1(\as2650.stack[12][7] ),
    .A2(_01811_),
    .B1(_02842_),
    .B2(\as2650.stack[13][7] ),
    .ZN(_02953_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08721_ (.A1(_02950_),
    .A2(_02952_),
    .A3(_02953_),
    .ZN(_02954_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08722_ (.A1(_02949_),
    .A2(_02954_),
    .ZN(_02955_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08723_ (.A1(\as2650.stack[0][7] ),
    .A2(_01811_),
    .B1(_02842_),
    .B2(\as2650.stack[1][7] ),
    .ZN(_02956_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08724_ (.I(_01962_),
    .Z(_02957_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08725_ (.A1(\as2650.stack[3][7] ),
    .A2(_02951_),
    .B1(_02957_),
    .B2(\as2650.stack[2][7] ),
    .ZN(_02958_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08726_ (.A1(_02834_),
    .A2(_02956_),
    .A3(_02958_),
    .ZN(_02959_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08727_ (.A1(\as2650.stack[7][7] ),
    .A2(_02951_),
    .B1(_02957_),
    .B2(\as2650.stack[6][7] ),
    .ZN(_02960_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08728_ (.I(_01810_),
    .Z(_02961_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08729_ (.I(_01953_),
    .Z(_02962_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08730_ (.A1(\as2650.stack[4][7] ),
    .A2(_02961_),
    .B1(_02962_),
    .B2(\as2650.stack[5][7] ),
    .ZN(_02963_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08731_ (.A1(_02950_),
    .A2(_02960_),
    .A3(_02963_),
    .ZN(_02964_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08732_ (.A1(_02959_),
    .A2(_02964_),
    .B(_02817_),
    .ZN(_02965_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08733_ (.A1(_02946_),
    .A2(_02955_),
    .B(_02965_),
    .ZN(_02966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08734_ (.A1(_02816_),
    .A2(_02966_),
    .ZN(_02967_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08735_ (.A1(_02778_),
    .A2(_02900_),
    .A3(_02945_),
    .A4(_02967_),
    .Z(_02968_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08736_ (.A1(_02895_),
    .A2(_02968_),
    .ZN(_00178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08737_ (.I(_02726_),
    .Z(_02969_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08738_ (.I(_02969_),
    .Z(_02970_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _08739_ (.A1(_02444_),
    .A2(_02395_),
    .Z(_02971_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08740_ (.I(_02971_),
    .Z(_02972_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08741_ (.A1(\as2650.stack[15][0] ),
    .A2(_02972_),
    .ZN(_02973_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08742_ (.I(_01839_),
    .Z(_02974_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08743_ (.A1(_02974_),
    .A2(_02733_),
    .B(_02735_),
    .ZN(_02975_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08744_ (.A1(_02630_),
    .A2(_02970_),
    .B1(_02973_),
    .B2(_02975_),
    .ZN(_00179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08745_ (.A1(\as2650.stack[15][1] ),
    .A2(_02972_),
    .ZN(_02976_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08746_ (.I(_01857_),
    .Z(_02977_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08747_ (.I(_02721_),
    .Z(_02978_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08748_ (.I(_02727_),
    .Z(_02979_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08749_ (.A1(_02977_),
    .A2(_02978_),
    .B(_02979_),
    .ZN(_02980_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08750_ (.A1(_02637_),
    .A2(_02970_),
    .B1(_02976_),
    .B2(_02980_),
    .ZN(_00180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08751_ (.A1(\as2650.stack[15][2] ),
    .A2(_02972_),
    .ZN(_02981_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08752_ (.I(_01869_),
    .Z(_02982_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08753_ (.A1(_02982_),
    .A2(_02978_),
    .B(_02979_),
    .ZN(_02983_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08754_ (.A1(_02642_),
    .A2(_02970_),
    .B1(_02981_),
    .B2(_02983_),
    .ZN(_00181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08755_ (.A1(\as2650.stack[15][3] ),
    .A2(_02972_),
    .ZN(_02984_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08756_ (.I(_01880_),
    .Z(_02985_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08757_ (.A1(_02985_),
    .A2(_02978_),
    .B(_02979_),
    .ZN(_02986_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08758_ (.A1(_02645_),
    .A2(_02970_),
    .B1(_02984_),
    .B2(_02986_),
    .ZN(_00182_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08759_ (.I(_02727_),
    .Z(_02987_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08760_ (.I(_02971_),
    .Z(_02988_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08761_ (.A1(\as2650.stack[15][4] ),
    .A2(_02988_),
    .ZN(_02989_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08762_ (.I(_01891_),
    .Z(_02990_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08763_ (.A1(_02990_),
    .A2(_02978_),
    .B(_02979_),
    .ZN(_02991_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08764_ (.A1(_02648_),
    .A2(_02987_),
    .B1(_02989_),
    .B2(_02991_),
    .ZN(_00183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08765_ (.A1(\as2650.stack[15][5] ),
    .A2(_02988_),
    .ZN(_02992_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08766_ (.I(_01905_),
    .Z(_02993_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08767_ (.A1(_02993_),
    .A2(_02724_),
    .B(_02969_),
    .ZN(_02994_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08768_ (.A1(_02653_),
    .A2(_02987_),
    .B1(_02992_),
    .B2(_02994_),
    .ZN(_00184_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08769_ (.A1(\as2650.stack[15][6] ),
    .A2(_02988_),
    .ZN(_02995_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08770_ (.I(_01915_),
    .Z(_02996_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08771_ (.A1(_02996_),
    .A2(_02724_),
    .B(_02969_),
    .ZN(_02997_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08772_ (.A1(_02656_),
    .A2(_02987_),
    .B1(_02995_),
    .B2(_02997_),
    .ZN(_00185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08773_ (.A1(\as2650.stack[15][7] ),
    .A2(_02988_),
    .ZN(_02998_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08774_ (.I(_01924_),
    .Z(_02999_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08775_ (.A1(_02999_),
    .A2(_02724_),
    .B(_02969_),
    .ZN(_03000_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08776_ (.A1(_02659_),
    .A2(_02987_),
    .B1(_02998_),
    .B2(_03000_),
    .ZN(_00186_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08777_ (.I(_02454_),
    .Z(_03001_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08778_ (.I(_03001_),
    .Z(_03002_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08779_ (.A1(_02250_),
    .A2(_01938_),
    .ZN(_03003_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08780_ (.I(_03003_),
    .Z(_03004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08781_ (.A1(\as2650.stack[8][0] ),
    .A2(_03004_),
    .ZN(_03005_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _08782_ (.A1(_02974_),
    .A2(_02461_),
    .B(_02463_),
    .ZN(_03006_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08783_ (.A1(_02630_),
    .A2(_03002_),
    .B1(_03005_),
    .B2(_03006_),
    .ZN(_00187_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08784_ (.A1(\as2650.stack[8][1] ),
    .A2(_03004_),
    .ZN(_03007_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08785_ (.I(_02446_),
    .Z(_03008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08786_ (.I(_02455_),
    .Z(_03009_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08787_ (.A1(_02977_),
    .A2(_03008_),
    .B(_03009_),
    .ZN(_03010_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08788_ (.A1(_02637_),
    .A2(_03002_),
    .B1(_03007_),
    .B2(_03010_),
    .ZN(_00188_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08789_ (.A1(\as2650.stack[8][2] ),
    .A2(_03004_),
    .ZN(_03011_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08790_ (.A1(_02982_),
    .A2(_03008_),
    .B(_03009_),
    .ZN(_03012_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08791_ (.A1(_02642_),
    .A2(_03002_),
    .B1(_03011_),
    .B2(_03012_),
    .ZN(_00189_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08792_ (.A1(\as2650.stack[8][3] ),
    .A2(_03004_),
    .ZN(_03013_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08793_ (.A1(_02985_),
    .A2(_03008_),
    .B(_03009_),
    .ZN(_03014_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08794_ (.A1(_02645_),
    .A2(_03002_),
    .B1(_03013_),
    .B2(_03014_),
    .ZN(_00190_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08795_ (.I(_02455_),
    .Z(_03015_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08796_ (.I(_03003_),
    .Z(_03016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08797_ (.A1(\as2650.stack[8][4] ),
    .A2(_03016_),
    .ZN(_03017_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08798_ (.A1(_02990_),
    .A2(_03008_),
    .B(_03009_),
    .ZN(_03018_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08799_ (.A1(_02648_),
    .A2(_03015_),
    .B1(_03017_),
    .B2(_03018_),
    .ZN(_00191_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08800_ (.A1(\as2650.stack[8][5] ),
    .A2(_03016_),
    .ZN(_03019_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08801_ (.A1(_02993_),
    .A2(_02449_),
    .B(_03001_),
    .ZN(_03020_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08802_ (.A1(_02653_),
    .A2(_03015_),
    .B1(_03019_),
    .B2(_03020_),
    .ZN(_00192_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08803_ (.A1(\as2650.stack[8][6] ),
    .A2(_03016_),
    .ZN(_03021_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08804_ (.A1(_02996_),
    .A2(_02449_),
    .B(_03001_),
    .ZN(_03022_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08805_ (.A1(_02656_),
    .A2(_03015_),
    .B1(_03021_),
    .B2(_03022_),
    .ZN(_00193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08806_ (.A1(\as2650.stack[8][7] ),
    .A2(_03016_),
    .ZN(_03023_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08807_ (.A1(_02999_),
    .A2(_02449_),
    .B(_03001_),
    .ZN(_03024_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08808_ (.A1(_02659_),
    .A2(_03015_),
    .B1(_03023_),
    .B2(_03024_),
    .ZN(_00194_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08809_ (.I(_02319_),
    .Z(_03025_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08810_ (.I(_03025_),
    .Z(_03026_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08811_ (.I(_02394_),
    .Z(_03027_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08812_ (.A1(_02250_),
    .A2(_02253_),
    .A3(_03027_),
    .ZN(_03028_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08813_ (.I(_03028_),
    .Z(_03029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08814_ (.A1(\as2650.stack[11][0] ),
    .A2(_03029_),
    .ZN(_03030_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08815_ (.A1(_02974_),
    .A2(_02326_),
    .B(_02328_),
    .ZN(_03031_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08816_ (.A1(_02630_),
    .A2(_03026_),
    .B1(_03030_),
    .B2(_03031_),
    .ZN(_00195_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08817_ (.A1(\as2650.stack[11][1] ),
    .A2(_03029_),
    .ZN(_03032_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08818_ (.I(_02313_),
    .Z(_03033_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08819_ (.I(_02320_),
    .Z(_03034_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08820_ (.A1(_02977_),
    .A2(_03033_),
    .B(_03034_),
    .ZN(_03035_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08821_ (.A1(_02637_),
    .A2(_03026_),
    .B1(_03032_),
    .B2(_03035_),
    .ZN(_00196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08822_ (.A1(\as2650.stack[11][2] ),
    .A2(_03029_),
    .ZN(_03036_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08823_ (.A1(_02982_),
    .A2(_03033_),
    .B(_03034_),
    .ZN(_03037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08824_ (.A1(_02642_),
    .A2(_03026_),
    .B1(_03036_),
    .B2(_03037_),
    .ZN(_00197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08825_ (.A1(\as2650.stack[11][3] ),
    .A2(_03029_),
    .ZN(_03038_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08826_ (.A1(_02985_),
    .A2(_03033_),
    .B(_03034_),
    .ZN(_03039_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08827_ (.A1(_02645_),
    .A2(_03026_),
    .B1(_03038_),
    .B2(_03039_),
    .ZN(_00198_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08828_ (.I(_02320_),
    .Z(_03040_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08829_ (.I(_03028_),
    .Z(_03041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08830_ (.A1(\as2650.stack[11][4] ),
    .A2(_03041_),
    .ZN(_03042_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08831_ (.A1(_02990_),
    .A2(_03033_),
    .B(_03034_),
    .ZN(_03043_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08832_ (.A1(_02648_),
    .A2(_03040_),
    .B1(_03042_),
    .B2(_03043_),
    .ZN(_00199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08833_ (.A1(\as2650.stack[11][5] ),
    .A2(_03041_),
    .ZN(_03044_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08834_ (.A1(_02993_),
    .A2(_02316_),
    .B(_03025_),
    .ZN(_03045_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08835_ (.A1(_02653_),
    .A2(_03040_),
    .B1(_03044_),
    .B2(_03045_),
    .ZN(_00200_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08836_ (.A1(\as2650.stack[11][6] ),
    .A2(_03041_),
    .ZN(_03046_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08837_ (.A1(_02996_),
    .A2(_02316_),
    .B(_03025_),
    .ZN(_03047_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08838_ (.A1(_02656_),
    .A2(_03040_),
    .B1(_03046_),
    .B2(_03047_),
    .ZN(_00201_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08839_ (.A1(\as2650.stack[11][7] ),
    .A2(_03041_),
    .ZN(_03048_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08840_ (.A1(_02999_),
    .A2(_02316_),
    .B(_03025_),
    .ZN(_03049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08841_ (.A1(_02659_),
    .A2(_03040_),
    .B1(_03048_),
    .B2(_03049_),
    .ZN(_00202_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08842_ (.I(_01761_),
    .Z(_03050_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _08843_ (.I(_02709_),
    .Z(_03051_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08844_ (.I(_03051_),
    .Z(_03052_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08845_ (.A1(_02400_),
    .A2(_01816_),
    .A3(_02402_),
    .ZN(_03053_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08846_ (.I(_03053_),
    .Z(_03054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08847_ (.A1(\as2650.stack[1][0] ),
    .A2(_03054_),
    .ZN(_03055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _08848_ (.A1(_02974_),
    .A2(_02716_),
    .B(_02718_),
    .ZN(_03056_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08849_ (.A1(_03050_),
    .A2(_03052_),
    .B1(_03055_),
    .B2(_03056_),
    .ZN(_00203_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08850_ (.I(_01846_),
    .Z(_03057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08851_ (.A1(\as2650.stack[1][1] ),
    .A2(_03054_),
    .ZN(_03058_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08852_ (.I(_02704_),
    .Z(_03059_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08853_ (.I(_02710_),
    .Z(_03060_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08854_ (.A1(_02977_),
    .A2(_03059_),
    .B(_03060_),
    .ZN(_03061_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08855_ (.A1(_03057_),
    .A2(_03052_),
    .B1(_03058_),
    .B2(_03061_),
    .ZN(_00204_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08856_ (.I(_01862_),
    .Z(_03062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08857_ (.A1(\as2650.stack[1][2] ),
    .A2(_03054_),
    .ZN(_03063_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08858_ (.A1(_02982_),
    .A2(_03059_),
    .B(_03060_),
    .ZN(_03064_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08859_ (.A1(_03062_),
    .A2(_03052_),
    .B1(_03063_),
    .B2(_03064_),
    .ZN(_00205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08860_ (.I(_01873_),
    .Z(_03065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08861_ (.A1(\as2650.stack[1][3] ),
    .A2(_03054_),
    .ZN(_03066_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08862_ (.A1(_02985_),
    .A2(_03059_),
    .B(_03060_),
    .ZN(_03067_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08863_ (.A1(_03065_),
    .A2(_03052_),
    .B1(_03066_),
    .B2(_03067_),
    .ZN(_00206_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08864_ (.I(_01883_),
    .Z(_03068_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08865_ (.I(_02710_),
    .Z(_03069_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08866_ (.I(_03053_),
    .Z(_03070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08867_ (.A1(\as2650.stack[1][4] ),
    .A2(_03070_),
    .ZN(_03071_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08868_ (.A1(_02990_),
    .A2(_03059_),
    .B(_03060_),
    .ZN(_03072_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08869_ (.A1(_03068_),
    .A2(_03069_),
    .B1(_03071_),
    .B2(_03072_),
    .ZN(_00207_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08870_ (.I(_01895_),
    .Z(_03073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08871_ (.A1(\as2650.stack[1][5] ),
    .A2(_03070_),
    .ZN(_03074_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08872_ (.A1(_02993_),
    .A2(_02707_),
    .B(_03051_),
    .ZN(_03075_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08873_ (.A1(_03073_),
    .A2(_03069_),
    .B1(_03074_),
    .B2(_03075_),
    .ZN(_00208_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08874_ (.I(_01908_),
    .Z(_03076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08875_ (.A1(\as2650.stack[1][6] ),
    .A2(_03070_),
    .ZN(_03077_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08876_ (.A1(_02996_),
    .A2(_02707_),
    .B(_03051_),
    .ZN(_03078_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08877_ (.A1(_03076_),
    .A2(_03069_),
    .B1(_03077_),
    .B2(_03078_),
    .ZN(_00209_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08878_ (.I(_01918_),
    .Z(_03079_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08879_ (.A1(\as2650.stack[1][7] ),
    .A2(_03070_),
    .ZN(_03080_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08880_ (.A1(_02999_),
    .A2(_02707_),
    .B(_03051_),
    .ZN(_03081_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08881_ (.A1(_03079_),
    .A2(_03069_),
    .B1(_03080_),
    .B2(_03081_),
    .ZN(_00210_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08882_ (.A1(_05781_),
    .A2(_00901_),
    .ZN(_03082_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08883_ (.I(_03082_),
    .Z(_03083_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08884_ (.A1(_00814_),
    .A2(_01022_),
    .A3(_03083_),
    .ZN(_03084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08885_ (.I(_03084_),
    .Z(_03085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _08886_ (.A1(_01007_),
    .A2(_00475_),
    .ZN(_03086_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08887_ (.A1(_01060_),
    .A2(_03086_),
    .ZN(_03087_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08888_ (.A1(_00999_),
    .A2(_03087_),
    .ZN(_03088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08889_ (.I(_01038_),
    .Z(_03089_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _08890_ (.A1(_01034_),
    .A2(_03089_),
    .A3(_01056_),
    .A4(_03083_),
    .ZN(_03090_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _08891_ (.A1(_00622_),
    .A2(_01014_),
    .A3(_01017_),
    .ZN(_03091_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _08892_ (.A1(_01007_),
    .A2(_01763_),
    .A3(_03091_),
    .ZN(_03092_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _08893_ (.I(_03092_),
    .ZN(_03093_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _08894_ (.A1(_01028_),
    .A2(_01029_),
    .A3(_03083_),
    .Z(_03094_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08895_ (.I(_03094_),
    .Z(_03095_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _08896_ (.A1(_00673_),
    .A2(_01002_),
    .A3(_01004_),
    .A4(_03082_),
    .Z(_03096_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08897_ (.I(_03096_),
    .Z(_03097_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08898_ (.I(_03097_),
    .Z(_03098_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08899_ (.A1(_03093_),
    .A2(_03095_),
    .A3(_03098_),
    .ZN(_03099_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _08900_ (.A1(_03085_),
    .A2(_03088_),
    .A3(_03090_),
    .A4(_03099_),
    .ZN(_03100_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08901_ (.I(_03100_),
    .Z(_03101_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08902_ (.A1(_00989_),
    .A2(_03101_),
    .ZN(_03102_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08903_ (.I(_03102_),
    .Z(_03103_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08904_ (.I(_03095_),
    .Z(_03104_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08905_ (.I(_03090_),
    .Z(_03105_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08906_ (.I(_03084_),
    .Z(_03106_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _08907_ (.A1(_00671_),
    .A2(_01060_),
    .A3(_03086_),
    .ZN(_03107_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08908_ (.I(_03107_),
    .Z(_03108_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _08909_ (.I(_01079_),
    .Z(_03109_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08910_ (.I(_03107_),
    .Z(_03110_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08911_ (.I(_03096_),
    .Z(_03111_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08912_ (.A1(_00455_),
    .A2(_03111_),
    .ZN(_03112_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08913_ (.A1(_03109_),
    .A2(_03098_),
    .B(_03110_),
    .C(_03112_),
    .ZN(_03113_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _08914_ (.A1(_01060_),
    .A2(_01062_),
    .A3(_03086_),
    .ZN(_03114_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08915_ (.I(_03114_),
    .Z(_03115_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08916_ (.A1(_01072_),
    .A2(_03108_),
    .B(_03113_),
    .C(_03115_),
    .ZN(_03116_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08917_ (.I(_03084_),
    .Z(_03117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08918_ (.A1(_01070_),
    .A2(_03115_),
    .ZN(_03118_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08919_ (.A1(_03117_),
    .A2(_03118_),
    .ZN(_03119_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08920_ (.A1(_01054_),
    .A2(_03106_),
    .B1(_03116_),
    .B2(_03119_),
    .ZN(_03120_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08921_ (.I(_03090_),
    .Z(_03121_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _08922_ (.I(_03094_),
    .ZN(_03122_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08923_ (.A1(_01094_),
    .A2(_03121_),
    .B(_03122_),
    .ZN(_03123_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08924_ (.A1(_03105_),
    .A2(_03120_),
    .B(_03123_),
    .ZN(_03124_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08925_ (.A1(_01051_),
    .A2(_03104_),
    .B(_03124_),
    .ZN(_03125_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08926_ (.I(_03092_),
    .Z(_03126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08927_ (.I(_03126_),
    .Z(_03127_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08928_ (.I0(net82),
    .I1(_03125_),
    .S(_03127_),
    .Z(_03128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08929_ (.A1(_01008_),
    .A2(_01148_),
    .ZN(_03129_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _08930_ (.A1(_00978_),
    .A2(_03129_),
    .ZN(_03130_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _08931_ (.A1(_00989_),
    .A2(_03100_),
    .B(_03130_),
    .C(_00599_),
    .ZN(_03131_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08932_ (.I(_03131_),
    .Z(_03132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08933_ (.A1(\as2650.r123_2[1][0] ),
    .A2(_03132_),
    .ZN(_03133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08934_ (.I(_03130_),
    .Z(_03134_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08935_ (.I(_03134_),
    .Z(_03135_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08936_ (.A1(_01142_),
    .A2(_01146_),
    .A3(_03135_),
    .ZN(_03136_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08937_ (.A1(_03103_),
    .A2(_03128_),
    .B(_03133_),
    .C(_03136_),
    .ZN(_00211_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08938_ (.I(_03102_),
    .Z(_03137_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08939_ (.I(_03122_),
    .Z(_03138_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _08940_ (.A1(_01032_),
    .A2(_01039_),
    .A3(_03086_),
    .ZN(_03139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08941_ (.I(_03084_),
    .Z(_03140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08942_ (.I(_03107_),
    .Z(_03141_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08943_ (.A1(_00454_),
    .A2(_03111_),
    .ZN(_03142_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08944_ (.A1(_01216_),
    .A2(_03098_),
    .B(_03110_),
    .C(_03142_),
    .ZN(_03143_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08945_ (.I(_03114_),
    .Z(_03144_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08946_ (.A1(_01212_),
    .A2(_03141_),
    .B(_03143_),
    .C(_03144_),
    .ZN(_03145_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _08947_ (.A1(_00953_),
    .A2(_01061_),
    .A3(_03087_),
    .ZN(_03146_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08948_ (.I(_03146_),
    .Z(_03147_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08949_ (.A1(_01224_),
    .A2(_03147_),
    .B(_03085_),
    .ZN(_03148_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _08950_ (.A1(_01209_),
    .A2(_03140_),
    .B1(_03145_),
    .B2(_03148_),
    .ZN(_03149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08951_ (.A1(_01206_),
    .A2(_03139_),
    .ZN(_03150_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08952_ (.A1(_03139_),
    .A2(_03149_),
    .B(_03150_),
    .C(_03138_),
    .ZN(_03151_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08953_ (.A1(_01199_),
    .A2(_03138_),
    .B(_03151_),
    .ZN(_03152_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08954_ (.I0(net81),
    .I1(_03152_),
    .S(_03127_),
    .Z(_03153_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08955_ (.A1(_01240_),
    .A2(_03135_),
    .B1(_03132_),
    .B2(\as2650.r123_2[1][1] ),
    .ZN(_03154_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08956_ (.A1(_03137_),
    .A2(_03153_),
    .B(_03154_),
    .ZN(_00212_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _08957_ (.I(_01072_),
    .Z(_03155_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _08958_ (.A1(_00657_),
    .A2(_01763_),
    .A3(_01004_),
    .A4(_03083_),
    .ZN(_03156_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08959_ (.I(_03156_),
    .Z(_03157_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08960_ (.A1(_00953_),
    .A2(_00670_),
    .A3(_03087_),
    .ZN(_03158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08961_ (.A1(_00450_),
    .A2(_03156_),
    .ZN(_03159_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _08962_ (.A1(_02859_),
    .A2(_03157_),
    .B(_03158_),
    .C(_03159_),
    .ZN(_03160_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08963_ (.A1(_00434_),
    .A2(_03110_),
    .B(_03115_),
    .ZN(_03161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08964_ (.A1(_03155_),
    .A2(_03144_),
    .B1(_03160_),
    .B2(_03161_),
    .ZN(_03162_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08965_ (.I0(_01272_),
    .I1(_03162_),
    .S(_03117_),
    .Z(_03163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08966_ (.A1(_03105_),
    .A2(_03163_),
    .ZN(_03164_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08967_ (.A1(_01260_),
    .A2(_03139_),
    .B(_03095_),
    .ZN(_03165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _08968_ (.A1(_01254_),
    .A2(_03104_),
    .B1(_03164_),
    .B2(_03165_),
    .ZN(_03166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08969_ (.A1(net80),
    .A2(_03093_),
    .ZN(_03167_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _08970_ (.A1(_03093_),
    .A2(_03166_),
    .B(_03167_),
    .ZN(_03168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _08971_ (.A1(_01318_),
    .A2(_03135_),
    .B1(_03132_),
    .B2(\as2650.r123_2[1][2] ),
    .ZN(_03169_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08972_ (.A1(_03137_),
    .A2(_03168_),
    .B(_03169_),
    .ZN(_00213_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08973_ (.A1(_00452_),
    .A2(_03097_),
    .ZN(_03170_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _08974_ (.A1(_02863_),
    .A2(_03111_),
    .B(_03110_),
    .C(_03170_),
    .ZN(_03171_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _08975_ (.A1(_02885_),
    .A2(_03108_),
    .B(_03171_),
    .C(_03115_),
    .ZN(_03172_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08976_ (.I(_03146_),
    .Z(_03173_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08977_ (.A1(_01212_),
    .A2(_03173_),
    .B(_03085_),
    .ZN(_03174_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _08978_ (.A1(_01325_),
    .A2(_03106_),
    .B1(_03172_),
    .B2(_03174_),
    .C(_03121_),
    .ZN(_03175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08979_ (.A1(_01323_),
    .A2(_03139_),
    .ZN(_03176_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08980_ (.I(_03095_),
    .Z(_03177_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08981_ (.A1(_03175_),
    .A2(_03176_),
    .B(_03177_),
    .ZN(_03178_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08982_ (.A1(_01343_),
    .A2(_03104_),
    .B(_03178_),
    .ZN(_03179_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _08983_ (.I0(_01373_),
    .I1(_03179_),
    .S(_03127_),
    .Z(_03180_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _08984_ (.A1(_01230_),
    .A2(_01399_),
    .A3(_01400_),
    .ZN(_03181_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08985_ (.A1(_01398_),
    .A2(_03181_),
    .ZN(_03182_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _08986_ (.A1(\as2650.r123_2[1][3] ),
    .A2(_03132_),
    .B(_03182_),
    .ZN(_03183_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08987_ (.A1(_03137_),
    .A2(_03180_),
    .B(_03183_),
    .ZN(_00214_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08988_ (.I(_03181_),
    .Z(_03184_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _08989_ (.I(_03131_),
    .Z(_03185_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08990_ (.A1(\as2650.r123_2[1][4] ),
    .A2(_03185_),
    .ZN(_03186_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08991_ (.A1(_01485_),
    .A2(_03184_),
    .B(_03186_),
    .ZN(_03187_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _08992_ (.I(_03126_),
    .Z(_03188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _08993_ (.I(_03090_),
    .Z(_03189_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _08994_ (.A1(_00437_),
    .A2(_03097_),
    .ZN(_03190_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _08995_ (.A1(_01426_),
    .A2(_03111_),
    .B(_03107_),
    .C(_03190_),
    .ZN(_03191_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08996_ (.A1(_00425_),
    .A2(_03158_),
    .B(_03173_),
    .ZN(_03192_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _08997_ (.A1(_01262_),
    .A2(_03173_),
    .B1(_03191_),
    .B2(_03192_),
    .C(_03085_),
    .ZN(_03193_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _08998_ (.A1(_01420_),
    .A2(_03106_),
    .B(_03193_),
    .ZN(_03194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _08999_ (.A1(_03121_),
    .A2(_03194_),
    .ZN(_03195_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09000_ (.A1(_01416_),
    .A2(_03189_),
    .B(_03138_),
    .C(_03195_),
    .ZN(_03196_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09001_ (.A1(_01413_),
    .A2(_03104_),
    .ZN(_03197_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09002_ (.A1(_03188_),
    .A2(_03196_),
    .A3(_03197_),
    .ZN(_03198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09003_ (.A1(_01461_),
    .A2(_03093_),
    .ZN(_03199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09004_ (.A1(_03198_),
    .A2(_03199_),
    .ZN(_03200_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09005_ (.A1(_03103_),
    .A2(_03200_),
    .ZN(_03201_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09006_ (.A1(_03187_),
    .A2(_03201_),
    .Z(_03202_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09007_ (.I(_03202_),
    .Z(_00215_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09008_ (.I(_01535_),
    .Z(_03203_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09009_ (.A1(_03203_),
    .A2(_03157_),
    .ZN(_03204_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _09010_ (.A1(_00428_),
    .A2(_03157_),
    .B(_03108_),
    .C(_03204_),
    .ZN(_03205_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _09011_ (.A1(_02884_),
    .A2(_03141_),
    .B(_03205_),
    .C(_03144_),
    .ZN(_03206_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09012_ (.A1(_02885_),
    .A2(_03147_),
    .B(_03106_),
    .ZN(_03207_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _09013_ (.A1(_02146_),
    .A2(_03140_),
    .B1(_03206_),
    .B2(_03207_),
    .ZN(_03208_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09014_ (.A1(_01531_),
    .A2(_03105_),
    .B(_03122_),
    .ZN(_03209_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09015_ (.A1(_03189_),
    .A2(_03208_),
    .B(_03209_),
    .ZN(_03210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09016_ (.A1(_01526_),
    .A2(_03177_),
    .ZN(_03211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09017_ (.A1(_03126_),
    .A2(_03211_),
    .ZN(_03212_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _09018_ (.A1(_01514_),
    .A2(_03188_),
    .B1(_03210_),
    .B2(_03212_),
    .ZN(_03213_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09019_ (.A1(_01578_),
    .A2(_03135_),
    .B1(_03185_),
    .B2(\as2650.r123_2[1][5] ),
    .ZN(_03214_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09020_ (.A1(_03137_),
    .A2(_03213_),
    .B(_03214_),
    .ZN(_00216_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09021_ (.A1(_00424_),
    .A2(_03157_),
    .Z(_03215_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _09022_ (.A1(_02852_),
    .A2(_03098_),
    .B(_03108_),
    .C(_03215_),
    .ZN(_03216_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _09023_ (.A1(_02896_),
    .A2(_03141_),
    .B(_03216_),
    .C(_03144_),
    .ZN(_03217_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09024_ (.A1(_01617_),
    .A2(_03147_),
    .B(_03117_),
    .ZN(_03218_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _09025_ (.A1(_01616_),
    .A2(_03140_),
    .B1(_03217_),
    .B2(_03218_),
    .ZN(_03219_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09026_ (.A1(_01631_),
    .A2(_03121_),
    .B(_03122_),
    .ZN(_03220_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09027_ (.A1(_03189_),
    .A2(_03219_),
    .B(_03220_),
    .ZN(_03221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09028_ (.A1(_01614_),
    .A2(_03177_),
    .ZN(_03222_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09029_ (.A1(_03126_),
    .A2(_03222_),
    .ZN(_03223_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _09030_ (.A1(_01606_),
    .A2(_03188_),
    .B1(_03221_),
    .B2(_03223_),
    .ZN(_03224_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09031_ (.A1(_01668_),
    .A2(_03134_),
    .B1(_03185_),
    .B2(\as2650.r123_2[1][6] ),
    .ZN(_03225_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09032_ (.A1(_03103_),
    .A2(_03224_),
    .B(_03225_),
    .ZN(_00217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09033_ (.A1(\as2650.r123_2[1][7] ),
    .A2(_03185_),
    .ZN(_03226_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09034_ (.A1(_01758_),
    .A2(_03184_),
    .B(_03226_),
    .ZN(_03227_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09035_ (.I(_01694_),
    .Z(_03228_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09036_ (.I0(_00421_),
    .I1(_00602_),
    .S(_03097_),
    .Z(_03229_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09037_ (.A1(_03141_),
    .A2(_03229_),
    .ZN(_03230_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09038_ (.A1(_02883_),
    .A2(_03158_),
    .B(_03173_),
    .ZN(_03231_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _09039_ (.A1(_02884_),
    .A2(_03147_),
    .B1(_03230_),
    .B2(_03231_),
    .C(_03117_),
    .ZN(_03232_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09040_ (.A1(_02782_),
    .A2(_03140_),
    .B(_03232_),
    .ZN(_03233_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09041_ (.A1(_01713_),
    .A2(_03105_),
    .B(_03138_),
    .ZN(_03234_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09042_ (.A1(_03189_),
    .A2(_03233_),
    .B(_03234_),
    .ZN(_03235_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09043_ (.A1(_01702_),
    .A2(_03177_),
    .ZN(_03236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09044_ (.A1(_03127_),
    .A2(_03236_),
    .ZN(_03237_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_4 _09045_ (.A1(_03228_),
    .A2(_03188_),
    .B1(_03235_),
    .B2(_03237_),
    .ZN(_03238_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09046_ (.A1(_03103_),
    .A2(_03238_),
    .ZN(_03239_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09047_ (.A1(_03227_),
    .A2(_03239_),
    .Z(_03240_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09048_ (.I(_03240_),
    .Z(_00218_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09049_ (.A1(_01930_),
    .A2(_00984_),
    .B(_03129_),
    .ZN(_03241_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09050_ (.A1(_03134_),
    .A2(_03241_),
    .ZN(_03242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09051_ (.I(_03242_),
    .Z(_03243_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09052_ (.A1(_01230_),
    .A2(_00942_),
    .A3(_01400_),
    .ZN(_03244_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09053_ (.I(_03244_),
    .Z(_03245_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09054_ (.A1(_01990_),
    .A2(_03245_),
    .ZN(_03246_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09055_ (.A1(_01930_),
    .A2(_03129_),
    .ZN(_03247_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09056_ (.I(_03247_),
    .Z(_03248_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09057_ (.A1(_01142_),
    .A2(_03248_),
    .ZN(_03249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09058_ (.A1(_05763_),
    .A2(_03101_),
    .ZN(_03250_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09059_ (.I(_03250_),
    .Z(_03251_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _09060_ (.A1(_03243_),
    .A2(_03246_),
    .A3(_03249_),
    .B1(_03251_),
    .B2(_03128_),
    .ZN(_03252_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09061_ (.A1(_05718_),
    .A2(_03241_),
    .ZN(_03253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09062_ (.A1(_03253_),
    .A2(_03250_),
    .ZN(_03254_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09063_ (.I(_03254_),
    .Z(_03255_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09064_ (.I0(\as2650.r123_2[0][0] ),
    .I1(_03252_),
    .S(_03255_),
    .Z(_03256_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09065_ (.I(_03256_),
    .Z(_00219_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09066_ (.A1(_02042_),
    .A2(_03245_),
    .ZN(_03257_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09067_ (.A1(_01850_),
    .A2(_03248_),
    .ZN(_03258_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _09068_ (.A1(_03243_),
    .A2(_03257_),
    .A3(_03258_),
    .B1(_03251_),
    .B2(_03153_),
    .ZN(_03259_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09069_ (.I0(\as2650.r123_2[0][1] ),
    .I1(_03259_),
    .S(_03255_),
    .Z(_03260_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09070_ (.I(_03260_),
    .Z(_00220_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09071_ (.A1(_02065_),
    .A2(_03245_),
    .ZN(_03261_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09072_ (.A1(_01865_),
    .A2(_03248_),
    .ZN(_03262_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _09073_ (.A1(_03243_),
    .A2(_03261_),
    .A3(_03262_),
    .B1(_03251_),
    .B2(_03168_),
    .ZN(_03263_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09074_ (.I0(\as2650.r123_2[0][2] ),
    .I1(_03263_),
    .S(_03255_),
    .Z(_03264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09075_ (.I(_03264_),
    .Z(_00221_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09076_ (.I(_03242_),
    .Z(_03265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09077_ (.I(_03244_),
    .Z(_03266_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09078_ (.A1(_02095_),
    .A2(_03266_),
    .ZN(_03267_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09079_ (.A1(_02097_),
    .A2(_03248_),
    .ZN(_03268_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09080_ (.I(_03250_),
    .Z(_03269_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _09081_ (.A1(_03265_),
    .A2(_03267_),
    .A3(_03268_),
    .B1(_03269_),
    .B2(_03180_),
    .ZN(_03270_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09082_ (.I0(\as2650.r123_2[0][3] ),
    .I1(_03270_),
    .S(_03255_),
    .Z(_03271_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09083_ (.I(_03271_),
    .Z(_00222_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09084_ (.A1(_02118_),
    .A2(_03266_),
    .ZN(_03272_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09085_ (.A1(_02120_),
    .A2(_03247_),
    .ZN(_03273_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _09086_ (.A1(_03265_),
    .A2(_03272_),
    .A3(_03273_),
    .B1(_03269_),
    .B2(_03200_),
    .ZN(_03274_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09087_ (.I(_03254_),
    .Z(_03275_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09088_ (.I0(\as2650.r123_2[0][4] ),
    .I1(_03274_),
    .S(_03275_),
    .Z(_03276_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09089_ (.I(_03276_),
    .Z(_00223_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09090_ (.A1(_02144_),
    .A2(_03266_),
    .ZN(_03277_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09091_ (.A1(_02146_),
    .A2(_03247_),
    .ZN(_03278_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _09092_ (.A1(_03265_),
    .A2(_03277_),
    .A3(_03278_),
    .B1(_03269_),
    .B2(_03213_),
    .ZN(_03279_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09093_ (.I0(\as2650.r123_2[0][5] ),
    .I1(_03279_),
    .S(_03275_),
    .Z(_03280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09094_ (.I(_03280_),
    .Z(_00224_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09095_ (.A1(_02164_),
    .A2(_03266_),
    .ZN(_03281_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09096_ (.A1(_01616_),
    .A2(_03247_),
    .ZN(_03282_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _09097_ (.A1(_03265_),
    .A2(_03281_),
    .A3(_03282_),
    .B1(_03269_),
    .B2(_03224_),
    .ZN(_03283_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09098_ (.I0(\as2650.r123_2[0][6] ),
    .I1(_03283_),
    .S(_03275_),
    .Z(_03284_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09099_ (.I(_03284_),
    .Z(_00225_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09100_ (.I(_02782_),
    .Z(_03285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09101_ (.A1(_03285_),
    .A2(_03245_),
    .ZN(_03286_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09102_ (.A1(_03238_),
    .A2(_03251_),
    .B1(_03243_),
    .B2(_03286_),
    .ZN(_03287_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09103_ (.I0(\as2650.r123_2[0][7] ),
    .I1(_03287_),
    .S(_03275_),
    .Z(_03288_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09104_ (.I(_03288_),
    .Z(_00226_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09105_ (.I(_02472_),
    .Z(_03289_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09106_ (.I(_03289_),
    .Z(_03290_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09107_ (.A1(_02406_),
    .A2(_01784_),
    .ZN(_03291_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09108_ (.A1(_02250_),
    .A2(_03027_),
    .A3(_03291_),
    .ZN(_03292_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09109_ (.I(_03292_),
    .Z(_03293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09110_ (.A1(\as2650.stack[7][0] ),
    .A2(_03293_),
    .ZN(_03294_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09111_ (.I(_01839_),
    .Z(_03295_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09112_ (.A1(_03295_),
    .A2(_02479_),
    .B(_02481_),
    .ZN(_03296_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09113_ (.A1(_03050_),
    .A2(_03290_),
    .B1(_03294_),
    .B2(_03296_),
    .ZN(_00227_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09114_ (.A1(\as2650.stack[7][1] ),
    .A2(_03293_),
    .ZN(_03297_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09115_ (.I(_01857_),
    .Z(_03298_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09116_ (.I(_02467_),
    .Z(_03299_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09117_ (.I(_02473_),
    .Z(_03300_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09118_ (.A1(_03298_),
    .A2(_03299_),
    .B(_03300_),
    .ZN(_03301_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09119_ (.A1(_03057_),
    .A2(_03290_),
    .B1(_03297_),
    .B2(_03301_),
    .ZN(_00228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09120_ (.A1(\as2650.stack[7][2] ),
    .A2(_03293_),
    .ZN(_03302_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09121_ (.I(_01869_),
    .Z(_03303_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09122_ (.A1(_03303_),
    .A2(_03299_),
    .B(_03300_),
    .ZN(_03304_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09123_ (.A1(_03062_),
    .A2(_03290_),
    .B1(_03302_),
    .B2(_03304_),
    .ZN(_00229_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09124_ (.A1(\as2650.stack[7][3] ),
    .A2(_03293_),
    .ZN(_03305_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09125_ (.I(_01880_),
    .Z(_03306_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09126_ (.A1(_03306_),
    .A2(_03299_),
    .B(_03300_),
    .ZN(_03307_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09127_ (.A1(_03065_),
    .A2(_03290_),
    .B1(_03305_),
    .B2(_03307_),
    .ZN(_00230_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09128_ (.I(_02473_),
    .Z(_03308_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09129_ (.I(_03292_),
    .Z(_03309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09130_ (.A1(\as2650.stack[7][4] ),
    .A2(_03309_),
    .ZN(_03310_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09131_ (.I(_01891_),
    .Z(_03311_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09132_ (.A1(_03311_),
    .A2(_03299_),
    .B(_03300_),
    .ZN(_03312_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09133_ (.A1(_03068_),
    .A2(_03308_),
    .B1(_03310_),
    .B2(_03312_),
    .ZN(_00231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09134_ (.A1(\as2650.stack[7][5] ),
    .A2(_03309_),
    .ZN(_03313_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09135_ (.I(_01905_),
    .Z(_03314_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09136_ (.A1(_03314_),
    .A2(_02470_),
    .B(_03289_),
    .ZN(_03315_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09137_ (.A1(_03073_),
    .A2(_03308_),
    .B1(_03313_),
    .B2(_03315_),
    .ZN(_00232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09138_ (.A1(\as2650.stack[7][6] ),
    .A2(_03309_),
    .ZN(_03316_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09139_ (.I(_01915_),
    .Z(_03317_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09140_ (.A1(_03317_),
    .A2(_02470_),
    .B(_03289_),
    .ZN(_03318_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09141_ (.A1(_03076_),
    .A2(_03308_),
    .B1(_03316_),
    .B2(_03318_),
    .ZN(_00233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09142_ (.A1(\as2650.stack[7][7] ),
    .A2(_03309_),
    .ZN(_03319_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09143_ (.I(_01924_),
    .Z(_03320_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09144_ (.A1(_03320_),
    .A2(_02470_),
    .B(_03289_),
    .ZN(_03321_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09145_ (.A1(_03079_),
    .A2(_03308_),
    .B1(_03319_),
    .B2(_03321_),
    .ZN(_00234_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09146_ (.I(_03184_),
    .Z(_03322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09147_ (.A1(_01723_),
    .A2(_01756_),
    .ZN(_03323_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09148_ (.A1(_01720_),
    .A2(_01757_),
    .B(_03323_),
    .ZN(_03324_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09149_ (.A1(_01729_),
    .A2(_01754_),
    .Z(_03325_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09150_ (.A1(_01726_),
    .A2(_01755_),
    .B(_03325_),
    .ZN(_03326_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09151_ (.A1(_01732_),
    .A2(_01734_),
    .Z(_03327_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09152_ (.A1(_01735_),
    .A2(_01736_),
    .B(_03327_),
    .ZN(_03328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09153_ (.A1(_01737_),
    .A2(_01753_),
    .ZN(_03329_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09154_ (.A1(_01741_),
    .A2(_01752_),
    .B(_03329_),
    .ZN(_03330_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09155_ (.A1(_01660_),
    .A2(_01750_),
    .ZN(_03331_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09156_ (.A1(_01746_),
    .A2(_01751_),
    .ZN(_03332_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09157_ (.A1(_03331_),
    .A2(_03332_),
    .ZN(_03333_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09158_ (.A1(_05816_),
    .A2(_01742_),
    .B1(_01236_),
    .B2(_05757_),
    .ZN(_03334_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09159_ (.A1(_05757_),
    .A2(_05816_),
    .A3(_01742_),
    .A4(_01236_),
    .Z(_03335_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09160_ (.A1(_03334_),
    .A2(_03335_),
    .Z(_03336_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09161_ (.A1(_01748_),
    .A2(_01749_),
    .Z(_03337_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09162_ (.A1(_01748_),
    .A2(_01749_),
    .Z(_03338_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09163_ (.A1(_01747_),
    .A2(_03337_),
    .B(_03338_),
    .ZN(_03339_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09164_ (.A1(_05786_),
    .A2(_01383_),
    .A3(_05765_),
    .A4(_01389_),
    .Z(_03340_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09165_ (.A1(_01383_),
    .A2(_05766_),
    .B1(_01385_),
    .B2(_05786_),
    .ZN(_03341_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09166_ (.A1(_03340_),
    .A2(_03341_),
    .Z(_03342_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09167_ (.A1(_05854_),
    .A2(_01311_),
    .ZN(_03343_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09168_ (.A1(_03342_),
    .A2(_03343_),
    .ZN(_03344_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09169_ (.A1(_03336_),
    .A2(_03339_),
    .A3(_03344_),
    .ZN(_03345_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09170_ (.I(_03345_),
    .ZN(_03346_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09171_ (.A1(_03333_),
    .A2(_03346_),
    .Z(_03347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09172_ (.A1(_01744_),
    .A2(_01745_),
    .ZN(_03348_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09173_ (.A1(_01744_),
    .A2(_01745_),
    .ZN(_03349_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09174_ (.A1(_01743_),
    .A2(_03348_),
    .B(_03349_),
    .ZN(_03350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09175_ (.A1(_05808_),
    .A2(_01733_),
    .ZN(_03351_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09176_ (.A1(_03350_),
    .A2(_03351_),
    .ZN(_03352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09177_ (.A1(_05797_),
    .A2(_01468_),
    .ZN(_03353_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09178_ (.A1(_03352_),
    .A2(_03353_),
    .ZN(_03354_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09179_ (.A1(_03347_),
    .A2(_03354_),
    .Z(_03355_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09180_ (.A1(_03330_),
    .A2(_03355_),
    .Z(_03356_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09181_ (.A1(_03328_),
    .A2(_03356_),
    .ZN(_03357_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09182_ (.A1(_03326_),
    .A2(_03357_),
    .Z(_03358_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _09183_ (.A1(_03324_),
    .A2(_03358_),
    .ZN(_03359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09184_ (.A1(_00947_),
    .A2(_03101_),
    .ZN(_03360_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09185_ (.I(_03360_),
    .Z(_03361_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _09186_ (.A1(_00947_),
    .A2(_03101_),
    .B(_03134_),
    .C(_00909_),
    .ZN(_03362_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09187_ (.I(_03362_),
    .Z(_03363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09188_ (.A1(\as2650.r123_2[2][0] ),
    .A2(_03363_),
    .ZN(_03364_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _09189_ (.A1(_03322_),
    .A2(_03359_),
    .B1(_03361_),
    .B2(_03128_),
    .C(_03364_),
    .ZN(_00235_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09190_ (.I(_03360_),
    .Z(_03365_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09191_ (.A1(_03326_),
    .A2(_03357_),
    .ZN(_03366_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09192_ (.A1(_03324_),
    .A2(_03358_),
    .B(_03366_),
    .ZN(_03367_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09193_ (.A1(_03330_),
    .A2(_03355_),
    .ZN(_03368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09194_ (.A1(_03328_),
    .A2(_03356_),
    .ZN(_03369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09195_ (.A1(_03368_),
    .A2(_03369_),
    .ZN(_03370_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09196_ (.A1(_03350_),
    .A2(_03351_),
    .Z(_03371_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09197_ (.A1(_03352_),
    .A2(_03353_),
    .B(_03371_),
    .ZN(_03372_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09198_ (.A1(_03333_),
    .A2(_03345_),
    .Z(_03373_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09199_ (.A1(_03347_),
    .A2(_03354_),
    .B(_03373_),
    .ZN(_03374_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09200_ (.I(_03344_),
    .ZN(_03375_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09201_ (.A1(_03339_),
    .A2(_03375_),
    .ZN(_03376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09202_ (.A1(_03339_),
    .A2(_03375_),
    .ZN(_03377_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09203_ (.A1(_03336_),
    .A2(_03376_),
    .B(_03377_),
    .ZN(_03378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09204_ (.A1(_05808_),
    .A2(_02228_),
    .ZN(_03379_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09205_ (.A1(_03342_),
    .A2(_03343_),
    .ZN(_03380_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09206_ (.A1(_03340_),
    .A2(_03380_),
    .ZN(_03381_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09207_ (.A1(\as2650.r0[6] ),
    .A2(\as2650.r0[2] ),
    .A3(_05765_),
    .A4(_01389_),
    .Z(_03382_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09208_ (.A1(_05815_),
    .A2(_05766_),
    .B1(_01389_),
    .B2(\as2650.r0[6] ),
    .ZN(_03383_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09209_ (.A1(_03382_),
    .A2(_03383_),
    .Z(_03384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09210_ (.A1(\as2650.r0[7] ),
    .A2(_01386_),
    .ZN(_03385_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09211_ (.A1(_03384_),
    .A2(_03385_),
    .ZN(_03386_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09212_ (.A1(_03381_),
    .A2(_03386_),
    .Z(_03387_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09213_ (.A1(_03379_),
    .A2(_03387_),
    .ZN(_03388_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09214_ (.A1(_03378_),
    .A2(_03388_),
    .Z(_03389_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09215_ (.A1(_01418_),
    .A2(_01733_),
    .ZN(_03390_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09216_ (.A1(_05787_),
    .A2(_01640_),
    .ZN(_03391_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09217_ (.A1(_03335_),
    .A2(_03390_),
    .A3(_03391_),
    .Z(_03392_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09218_ (.A1(_03389_),
    .A2(_03392_),
    .Z(_03393_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09219_ (.A1(_03374_),
    .A2(_03393_),
    .Z(_03394_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09220_ (.A1(_03372_),
    .A2(_03394_),
    .Z(_03395_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09221_ (.A1(_03370_),
    .A2(_03395_),
    .ZN(_03396_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _09222_ (.A1(_03367_),
    .A2(_03396_),
    .ZN(_03397_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09223_ (.I(_03184_),
    .Z(_03398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09224_ (.A1(\as2650.r123_2[2][1] ),
    .A2(_03363_),
    .ZN(_03399_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _09225_ (.A1(_03153_),
    .A2(_03365_),
    .B1(_03397_),
    .B2(_03398_),
    .C(_03399_),
    .ZN(_00236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09226_ (.A1(_03370_),
    .A2(_03395_),
    .ZN(_03400_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09227_ (.A1(_03367_),
    .A2(_03396_),
    .B(_03400_),
    .ZN(_03401_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09228_ (.A1(_03374_),
    .A2(_03393_),
    .Z(_03402_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09229_ (.A1(_03372_),
    .A2(_03394_),
    .B(_03402_),
    .ZN(_03403_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09230_ (.A1(_01419_),
    .A2(_02223_),
    .B(_03335_),
    .ZN(_03404_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09231_ (.A1(_01420_),
    .A2(_02223_),
    .A3(_03335_),
    .ZN(_03405_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09232_ (.A1(_03404_),
    .A2(_03391_),
    .B(_03405_),
    .ZN(_03406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09233_ (.A1(_03378_),
    .A2(_03388_),
    .ZN(_03407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09234_ (.A1(_03389_),
    .A2(_03392_),
    .ZN(_03408_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09235_ (.A1(_03407_),
    .A2(_03408_),
    .ZN(_03409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09236_ (.A1(_05855_),
    .A2(_01640_),
    .ZN(_03410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09237_ (.A1(_01493_),
    .A2(_02222_),
    .ZN(_03411_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09238_ (.A1(_03410_),
    .A2(_03411_),
    .ZN(_03412_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09239_ (.A1(_03410_),
    .A2(_03411_),
    .Z(_03413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09240_ (.A1(_03412_),
    .A2(_03413_),
    .ZN(_03414_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09241_ (.A1(_05809_),
    .A2(_02228_),
    .A3(_03387_),
    .ZN(_03415_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09242_ (.A1(_03381_),
    .A2(_03386_),
    .B(_03415_),
    .ZN(_03416_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09243_ (.A1(_05807_),
    .A2(_05766_),
    .ZN(_03417_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09244_ (.A1(_05758_),
    .A2(_01476_),
    .ZN(_03418_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09245_ (.A1(_03384_),
    .A2(_03385_),
    .ZN(_03419_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09246_ (.A1(_03382_),
    .A2(_03419_),
    .ZN(_03420_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09247_ (.A1(_03417_),
    .A2(_03418_),
    .A3(_03420_),
    .ZN(_03421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09248_ (.A1(_05797_),
    .A2(_02228_),
    .ZN(_03422_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09249_ (.A1(_03421_),
    .A2(_03422_),
    .ZN(_03423_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09250_ (.A1(_03416_),
    .A2(_03423_),
    .ZN(_03424_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09251_ (.A1(_03414_),
    .A2(_03424_),
    .Z(_03425_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09252_ (.A1(_03409_),
    .A2(_03425_),
    .Z(_03426_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09253_ (.A1(_03406_),
    .A2(_03426_),
    .ZN(_03427_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09254_ (.A1(_03403_),
    .A2(_03427_),
    .Z(_03428_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _09255_ (.A1(_03401_),
    .A2(_03428_),
    .ZN(_03429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09256_ (.A1(\as2650.r123_2[2][2] ),
    .A2(_03363_),
    .ZN(_03430_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _09257_ (.A1(_03168_),
    .A2(_03365_),
    .B1(_03429_),
    .B2(_03398_),
    .C(_03430_),
    .ZN(_00237_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09258_ (.A1(_03403_),
    .A2(_03427_),
    .ZN(_03431_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09259_ (.A1(_03401_),
    .A2(_03428_),
    .B(_03431_),
    .ZN(_03432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09260_ (.A1(_03409_),
    .A2(_03425_),
    .ZN(_03433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09261_ (.A1(_03406_),
    .A2(_03426_),
    .ZN(_03434_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09262_ (.A1(_03416_),
    .A2(_03423_),
    .ZN(_03435_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09263_ (.A1(_03414_),
    .A2(_03424_),
    .B(_03435_),
    .ZN(_03436_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09264_ (.A1(_05758_),
    .A2(_01724_),
    .ZN(_03437_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09265_ (.A1(_01587_),
    .A2(_02222_),
    .ZN(_03438_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09266_ (.A1(_03437_),
    .A2(_03438_),
    .ZN(_03439_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _09267_ (.A1(_03437_),
    .A2(_03438_),
    .Z(_03440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09268_ (.A1(_03439_),
    .A2(_03440_),
    .ZN(_03441_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09269_ (.A1(_03417_),
    .A2(_03418_),
    .ZN(_03442_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09270_ (.A1(_03417_),
    .A2(_03418_),
    .Z(_03443_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09271_ (.A1(_01419_),
    .A2(_02229_),
    .A3(_03421_),
    .ZN(_03444_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _09272_ (.A1(_03442_),
    .A2(_03443_),
    .A3(_03420_),
    .B(_03444_),
    .ZN(_03445_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09273_ (.A1(_01418_),
    .A2(_05767_),
    .Z(_03446_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09274_ (.A1(_01418_),
    .A2(_03442_),
    .ZN(_03447_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09275_ (.A1(_03442_),
    .A2(_03446_),
    .B(_03447_),
    .ZN(_03448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09276_ (.A1(_05787_),
    .A2(_02229_),
    .ZN(_03449_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09277_ (.A1(_03448_),
    .A2(_03449_),
    .ZN(_03450_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09278_ (.A1(_03445_),
    .A2(_03450_),
    .Z(_03451_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09279_ (.A1(_03441_),
    .A2(_03451_),
    .Z(_03452_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09280_ (.A1(_03436_),
    .A2(_03452_),
    .Z(_03453_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09281_ (.A1(_03413_),
    .A2(_03453_),
    .Z(_03454_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09282_ (.A1(_03433_),
    .A2(_03434_),
    .B(_03454_),
    .ZN(_03455_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _09283_ (.A1(_03433_),
    .A2(_03434_),
    .A3(_03454_),
    .Z(_03456_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09284_ (.A1(_03455_),
    .A2(_03456_),
    .ZN(_03457_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _09285_ (.A1(_03432_),
    .A2(_03457_),
    .Z(_03458_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09286_ (.A1(\as2650.r123_2[2][3] ),
    .A2(_03363_),
    .ZN(_03459_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _09287_ (.A1(_03180_),
    .A2(_03365_),
    .B1(_03458_),
    .B2(_03398_),
    .C(_03459_),
    .ZN(_00238_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09288_ (.I(_03455_),
    .ZN(_03460_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09289_ (.A1(_03432_),
    .A2(_03456_),
    .B(_03460_),
    .ZN(_03461_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09290_ (.I(_03453_),
    .ZN(_03462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09291_ (.A1(_03436_),
    .A2(_03452_),
    .ZN(_03463_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09292_ (.A1(_03413_),
    .A2(_03462_),
    .B(_03463_),
    .ZN(_03464_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09293_ (.I(_03450_),
    .ZN(_03465_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09294_ (.A1(_03445_),
    .A2(_03465_),
    .ZN(_03466_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09295_ (.A1(_03441_),
    .A2(_03451_),
    .B(_03466_),
    .ZN(_03467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09296_ (.A1(_01673_),
    .A2(_02222_),
    .ZN(_03468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09297_ (.A1(_05855_),
    .A2(_02229_),
    .ZN(_03469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09298_ (.A1(_01493_),
    .A2(_05767_),
    .ZN(_03470_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09299_ (.A1(_03469_),
    .A2(_03470_),
    .Z(_03471_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09300_ (.A1(_03448_),
    .A2(_03449_),
    .B(_03447_),
    .ZN(_03472_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09301_ (.A1(_03468_),
    .A2(_03471_),
    .A3(_03472_),
    .ZN(_03473_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09302_ (.A1(_03467_),
    .A2(_03473_),
    .ZN(_03474_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09303_ (.A1(_03440_),
    .A2(_03474_),
    .Z(_03475_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09304_ (.A1(_03464_),
    .A2(_03475_),
    .Z(_03476_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09305_ (.A1(_03461_),
    .A2(_03476_),
    .ZN(_03477_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09306_ (.I(_03362_),
    .Z(_03478_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09307_ (.A1(\as2650.r123_2[2][4] ),
    .A2(_03478_),
    .ZN(_03479_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _09308_ (.A1(_03200_),
    .A2(_03365_),
    .B1(_03477_),
    .B2(_03398_),
    .C(_03479_),
    .ZN(_00239_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09309_ (.A1(_03464_),
    .A2(_03475_),
    .Z(_03480_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09310_ (.A1(_03461_),
    .A2(_03476_),
    .B(_03480_),
    .ZN(_03481_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09311_ (.A1(_03471_),
    .A2(_03472_),
    .ZN(_03482_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09312_ (.A1(_03471_),
    .A2(_03472_),
    .ZN(_03483_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09313_ (.A1(_03468_),
    .A2(_03482_),
    .B(_03483_),
    .ZN(_03484_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _09314_ (.A1(_03469_),
    .A2(_03470_),
    .Z(_03485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09315_ (.I(_05767_),
    .Z(_03486_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09316_ (.A1(_01615_),
    .A2(_03486_),
    .B1(_02230_),
    .B2(_01673_),
    .ZN(_03487_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09317_ (.A1(_01673_),
    .A2(_01587_),
    .A3(_03486_),
    .A4(_02230_),
    .Z(_03488_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09318_ (.A1(_03487_),
    .A2(_03488_),
    .B(_03485_),
    .ZN(_03489_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09319_ (.A1(_01674_),
    .A2(_03485_),
    .B(_03489_),
    .ZN(_03490_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09320_ (.A1(_03484_),
    .A2(_03490_),
    .ZN(_03491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09321_ (.A1(_03467_),
    .A2(_03473_),
    .ZN(_03492_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09322_ (.A1(_03440_),
    .A2(_03474_),
    .B(_03492_),
    .ZN(_03493_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09323_ (.A1(_03491_),
    .A2(_03493_),
    .ZN(_03494_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09324_ (.A1(_03481_),
    .A2(_03494_),
    .ZN(_03495_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09325_ (.A1(\as2650.r123_2[2][5] ),
    .A2(_03478_),
    .ZN(_03496_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _09326_ (.A1(_03213_),
    .A2(_03361_),
    .B1(_03495_),
    .B2(_03322_),
    .C(_03496_),
    .ZN(_00240_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _09327_ (.A1(_01703_),
    .A2(_03485_),
    .B(_03484_),
    .C(_03489_),
    .ZN(_03497_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09328_ (.A1(_03491_),
    .A2(_03493_),
    .ZN(_03498_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09329_ (.A1(_03481_),
    .A2(_03494_),
    .B(_03498_),
    .ZN(_03499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09330_ (.A1(_03486_),
    .A2(_03469_),
    .ZN(_03500_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09331_ (.I0(_03485_),
    .I1(_03500_),
    .S(_02782_),
    .Z(_03501_));
 gf180mcu_fd_sc_mcu7t5v0__xnor3_1 _09332_ (.A1(_03497_),
    .A2(_03499_),
    .A3(_03501_),
    .ZN(_03502_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09333_ (.A1(\as2650.r123_2[2][6] ),
    .A2(_03478_),
    .ZN(_03503_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _09334_ (.A1(_03224_),
    .A2(_03361_),
    .B1(_03502_),
    .B2(_03322_),
    .C(_03503_),
    .ZN(_00241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09335_ (.A1(_03497_),
    .A2(_03501_),
    .ZN(_03504_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09336_ (.A1(_03497_),
    .A2(_03501_),
    .ZN(_03505_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _09337_ (.A1(_03499_),
    .A2(_03504_),
    .B(_03505_),
    .C(_03488_),
    .ZN(_03506_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09338_ (.A1(\as2650.r123_2[2][7] ),
    .A2(_03478_),
    .ZN(_03507_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _09339_ (.A1(_03238_),
    .A2(_03361_),
    .B1(_03506_),
    .B2(_03322_),
    .C(_03507_),
    .ZN(_00242_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09340_ (.I(_02668_),
    .Z(_03508_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09341_ (.I(_03508_),
    .Z(_03509_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09342_ (.I(_01807_),
    .Z(_03510_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09343_ (.A1(_03510_),
    .A2(_03027_),
    .A3(_02402_),
    .ZN(_03511_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09344_ (.I(_03511_),
    .Z(_03512_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09345_ (.A1(\as2650.stack[3][0] ),
    .A2(_03512_),
    .ZN(_03513_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09346_ (.A1(_03295_),
    .A2(_02675_),
    .B(_02677_),
    .ZN(_03514_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09347_ (.A1(_03050_),
    .A2(_03509_),
    .B1(_03513_),
    .B2(_03514_),
    .ZN(_00243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09348_ (.A1(\as2650.stack[3][1] ),
    .A2(_03512_),
    .ZN(_03515_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09349_ (.I(_02662_),
    .Z(_03516_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09350_ (.I(_02669_),
    .Z(_03517_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09351_ (.A1(_03298_),
    .A2(_03516_),
    .B(_03517_),
    .ZN(_03518_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09352_ (.A1(_03057_),
    .A2(_03509_),
    .B1(_03515_),
    .B2(_03518_),
    .ZN(_00244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09353_ (.A1(\as2650.stack[3][2] ),
    .A2(_03512_),
    .ZN(_03519_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09354_ (.A1(_03303_),
    .A2(_03516_),
    .B(_03517_),
    .ZN(_03520_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09355_ (.A1(_03062_),
    .A2(_03509_),
    .B1(_03519_),
    .B2(_03520_),
    .ZN(_00245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09356_ (.A1(\as2650.stack[3][3] ),
    .A2(_03512_),
    .ZN(_03521_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09357_ (.A1(_03306_),
    .A2(_03516_),
    .B(_03517_),
    .ZN(_03522_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09358_ (.A1(_03065_),
    .A2(_03509_),
    .B1(_03521_),
    .B2(_03522_),
    .ZN(_00246_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09359_ (.I(_02669_),
    .Z(_03523_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09360_ (.I(_03511_),
    .Z(_03524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09361_ (.A1(\as2650.stack[3][4] ),
    .A2(_03524_),
    .ZN(_03525_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09362_ (.A1(_03311_),
    .A2(_03516_),
    .B(_03517_),
    .ZN(_03526_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09363_ (.A1(_03068_),
    .A2(_03523_),
    .B1(_03525_),
    .B2(_03526_),
    .ZN(_00247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09364_ (.A1(\as2650.stack[3][5] ),
    .A2(_03524_),
    .ZN(_03527_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09365_ (.A1(_03314_),
    .A2(_02665_),
    .B(_03508_),
    .ZN(_03528_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09366_ (.A1(_03073_),
    .A2(_03523_),
    .B1(_03527_),
    .B2(_03528_),
    .ZN(_00248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09367_ (.A1(\as2650.stack[3][6] ),
    .A2(_03524_),
    .ZN(_03529_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09368_ (.A1(_03317_),
    .A2(_02665_),
    .B(_03508_),
    .ZN(_03530_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09369_ (.A1(_03076_),
    .A2(_03523_),
    .B1(_03529_),
    .B2(_03530_),
    .ZN(_00249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09370_ (.A1(\as2650.stack[3][7] ),
    .A2(_03524_),
    .ZN(_03531_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09371_ (.A1(_03320_),
    .A2(_02665_),
    .B(_03508_),
    .ZN(_03532_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09372_ (.A1(_03079_),
    .A2(_03523_),
    .B1(_03531_),
    .B2(_03532_),
    .ZN(_00250_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09373_ (.I(_02600_),
    .Z(_03533_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09374_ (.I(_03533_),
    .Z(_03534_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09375_ (.A1(_03510_),
    .A2(_01816_),
    .A3(_03291_),
    .ZN(_03535_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09376_ (.I(_03535_),
    .Z(_03536_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09377_ (.A1(\as2650.stack[5][0] ),
    .A2(_03536_),
    .ZN(_03537_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09378_ (.A1(_03295_),
    .A2(_02607_),
    .B(_02609_),
    .ZN(_03538_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09379_ (.A1(_03050_),
    .A2(_03534_),
    .B1(_03537_),
    .B2(_03538_),
    .ZN(_00251_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09380_ (.A1(\as2650.stack[5][1] ),
    .A2(_03536_),
    .ZN(_03539_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09381_ (.I(_02595_),
    .Z(_03540_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09382_ (.I(_02601_),
    .Z(_03541_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09383_ (.A1(_03298_),
    .A2(_03540_),
    .B(_03541_),
    .ZN(_03542_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09384_ (.A1(_03057_),
    .A2(_03534_),
    .B1(_03539_),
    .B2(_03542_),
    .ZN(_00252_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09385_ (.A1(\as2650.stack[5][2] ),
    .A2(_03536_),
    .ZN(_03543_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09386_ (.A1(_03303_),
    .A2(_03540_),
    .B(_03541_),
    .ZN(_03544_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09387_ (.A1(_03062_),
    .A2(_03534_),
    .B1(_03543_),
    .B2(_03544_),
    .ZN(_00253_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09388_ (.A1(\as2650.stack[5][3] ),
    .A2(_03536_),
    .ZN(_03545_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09389_ (.A1(_03306_),
    .A2(_03540_),
    .B(_03541_),
    .ZN(_03546_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09390_ (.A1(_03065_),
    .A2(_03534_),
    .B1(_03545_),
    .B2(_03546_),
    .ZN(_00254_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09391_ (.I(_02601_),
    .Z(_03547_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09392_ (.I(_03535_),
    .Z(_03548_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09393_ (.A1(\as2650.stack[5][4] ),
    .A2(_03548_),
    .ZN(_03549_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09394_ (.A1(_03311_),
    .A2(_03540_),
    .B(_03541_),
    .ZN(_03550_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09395_ (.A1(_03068_),
    .A2(_03547_),
    .B1(_03549_),
    .B2(_03550_),
    .ZN(_00255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09396_ (.A1(\as2650.stack[5][5] ),
    .A2(_03548_),
    .ZN(_03551_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09397_ (.A1(_03314_),
    .A2(_02598_),
    .B(_03533_),
    .ZN(_03552_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09398_ (.A1(_03073_),
    .A2(_03547_),
    .B1(_03551_),
    .B2(_03552_),
    .ZN(_00256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09399_ (.A1(\as2650.stack[5][6] ),
    .A2(_03548_),
    .ZN(_03553_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09400_ (.A1(_03317_),
    .A2(_02598_),
    .B(_03533_),
    .ZN(_03554_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09401_ (.A1(_03076_),
    .A2(_03547_),
    .B1(_03553_),
    .B2(_03554_),
    .ZN(_00257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09402_ (.A1(\as2650.stack[5][7] ),
    .A2(_03548_),
    .ZN(_03555_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09403_ (.A1(_03320_),
    .A2(_02598_),
    .B(_03533_),
    .ZN(_03556_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09404_ (.A1(_03079_),
    .A2(_03547_),
    .B1(_03555_),
    .B2(_03556_),
    .ZN(_00258_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09405_ (.I(_01760_),
    .Z(_03557_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09406_ (.I(_02618_),
    .Z(_03558_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09407_ (.I(_03558_),
    .Z(_03559_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09408_ (.A1(_02399_),
    .A2(_02400_),
    .A3(_03291_),
    .ZN(_03560_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09409_ (.I(_03560_),
    .Z(_03561_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09410_ (.A1(\as2650.stack[4][0] ),
    .A2(_03561_),
    .ZN(_03562_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09411_ (.A1(_03295_),
    .A2(_02625_),
    .B(_02627_),
    .ZN(_03563_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09412_ (.A1(_03557_),
    .A2(_03559_),
    .B1(_03562_),
    .B2(_03563_),
    .ZN(_00259_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09413_ (.I(_01845_),
    .Z(_03564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09414_ (.A1(\as2650.stack[4][1] ),
    .A2(_03561_),
    .ZN(_03565_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09415_ (.I(_02612_),
    .Z(_03566_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09416_ (.I(_02619_),
    .Z(_03567_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09417_ (.A1(_03298_),
    .A2(_03566_),
    .B(_03567_),
    .ZN(_03568_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09418_ (.A1(_03564_),
    .A2(_03559_),
    .B1(_03565_),
    .B2(_03568_),
    .ZN(_00260_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09419_ (.I(_01861_),
    .Z(_03569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09420_ (.A1(\as2650.stack[4][2] ),
    .A2(_03561_),
    .ZN(_03570_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09421_ (.A1(_03303_),
    .A2(_03566_),
    .B(_03567_),
    .ZN(_03571_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09422_ (.A1(_03569_),
    .A2(_03559_),
    .B1(_03570_),
    .B2(_03571_),
    .ZN(_00261_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09423_ (.I(_01872_),
    .Z(_03572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09424_ (.A1(\as2650.stack[4][3] ),
    .A2(_03561_),
    .ZN(_03573_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09425_ (.A1(_03306_),
    .A2(_03566_),
    .B(_03567_),
    .ZN(_03574_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09426_ (.A1(_03572_),
    .A2(_03559_),
    .B1(_03573_),
    .B2(_03574_),
    .ZN(_00262_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09427_ (.I(_01883_),
    .Z(_03575_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09428_ (.I(_02619_),
    .Z(_03576_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09429_ (.I(_03560_),
    .Z(_03577_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09430_ (.A1(\as2650.stack[4][4] ),
    .A2(_03577_),
    .ZN(_03578_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09431_ (.A1(_03311_),
    .A2(_03566_),
    .B(_03567_),
    .ZN(_03579_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09432_ (.A1(_03575_),
    .A2(_03576_),
    .B1(_03578_),
    .B2(_03579_),
    .ZN(_00263_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09433_ (.I(_01894_),
    .Z(_03580_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09434_ (.A1(\as2650.stack[4][5] ),
    .A2(_03577_),
    .ZN(_03581_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09435_ (.A1(_03314_),
    .A2(_02615_),
    .B(_03558_),
    .ZN(_03582_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09436_ (.A1(_03580_),
    .A2(_03576_),
    .B1(_03581_),
    .B2(_03582_),
    .ZN(_00264_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09437_ (.I(_01908_),
    .Z(_03583_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09438_ (.A1(\as2650.stack[4][6] ),
    .A2(_03577_),
    .ZN(_03584_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09439_ (.A1(_03317_),
    .A2(_02615_),
    .B(_03558_),
    .ZN(_03585_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09440_ (.A1(_03583_),
    .A2(_03576_),
    .B1(_03584_),
    .B2(_03585_),
    .ZN(_00265_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09441_ (.I(_01918_),
    .Z(_03586_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09442_ (.A1(\as2650.stack[4][7] ),
    .A2(_03577_),
    .ZN(_03587_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09443_ (.A1(_03320_),
    .A2(_02615_),
    .B(_03558_),
    .ZN(_03588_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09444_ (.A1(_03586_),
    .A2(_03576_),
    .B1(_03587_),
    .B2(_03588_),
    .ZN(_00266_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09445_ (.I(_02577_),
    .Z(_03589_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09446_ (.I(_03589_),
    .Z(_03590_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09447_ (.A1(_03510_),
    .A2(_02255_),
    .A3(_03291_),
    .ZN(_03591_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09448_ (.I(_03591_),
    .Z(_03592_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09449_ (.A1(\as2650.stack[6][0] ),
    .A2(_03592_),
    .ZN(_03593_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09450_ (.A1(_01840_),
    .A2(_02588_),
    .B(_02590_),
    .ZN(_03594_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09451_ (.A1(_03557_),
    .A2(_03590_),
    .B1(_03593_),
    .B2(_03594_),
    .ZN(_00267_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09452_ (.A1(\as2650.stack[6][1] ),
    .A2(_03592_),
    .ZN(_03595_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09453_ (.I(_02572_),
    .Z(_03596_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09454_ (.I(_02578_),
    .Z(_03597_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09455_ (.A1(_01858_),
    .A2(_03596_),
    .B(_03597_),
    .ZN(_03598_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09456_ (.A1(_03564_),
    .A2(_03590_),
    .B1(_03595_),
    .B2(_03598_),
    .ZN(_00268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09457_ (.A1(\as2650.stack[6][2] ),
    .A2(_03592_),
    .ZN(_03599_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09458_ (.A1(_01870_),
    .A2(_03596_),
    .B(_03597_),
    .ZN(_03600_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09459_ (.A1(_03569_),
    .A2(_03590_),
    .B1(_03599_),
    .B2(_03600_),
    .ZN(_00269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09460_ (.A1(\as2650.stack[6][3] ),
    .A2(_03592_),
    .ZN(_03601_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09461_ (.A1(_01881_),
    .A2(_03596_),
    .B(_03597_),
    .ZN(_03602_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09462_ (.A1(_03572_),
    .A2(_03590_),
    .B1(_03601_),
    .B2(_03602_),
    .ZN(_00270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09463_ (.I(_02578_),
    .Z(_03603_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09464_ (.I(_03591_),
    .Z(_03604_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09465_ (.A1(\as2650.stack[6][4] ),
    .A2(_03604_),
    .ZN(_03605_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09466_ (.A1(_01892_),
    .A2(_03596_),
    .B(_03597_),
    .ZN(_03606_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09467_ (.A1(_03575_),
    .A2(_03603_),
    .B1(_03605_),
    .B2(_03606_),
    .ZN(_00271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09468_ (.A1(\as2650.stack[6][5] ),
    .A2(_03604_),
    .ZN(_03607_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09469_ (.A1(_01906_),
    .A2(_02575_),
    .B(_03589_),
    .ZN(_03608_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09470_ (.A1(_03580_),
    .A2(_03603_),
    .B1(_03607_),
    .B2(_03608_),
    .ZN(_00272_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09471_ (.A1(\as2650.stack[6][6] ),
    .A2(_03604_),
    .ZN(_03609_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09472_ (.A1(_01916_),
    .A2(_02575_),
    .B(_03589_),
    .ZN(_03610_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09473_ (.A1(_03583_),
    .A2(_03603_),
    .B1(_03609_),
    .B2(_03610_),
    .ZN(_00273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09474_ (.A1(\as2650.stack[6][7] ),
    .A2(_03604_),
    .ZN(_03611_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09475_ (.A1(_01925_),
    .A2(_02575_),
    .B(_03589_),
    .ZN(_03612_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09476_ (.A1(_03586_),
    .A2(_03603_),
    .B1(_03611_),
    .B2(_03612_),
    .ZN(_00274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09477_ (.A1(_02738_),
    .A2(_02535_),
    .ZN(_03613_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _09478_ (.A1(_00599_),
    .A2(_00956_),
    .A3(_00937_),
    .A4(_03613_),
    .ZN(_03614_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09479_ (.I(_03614_),
    .Z(_03615_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09480_ (.I(_03615_),
    .Z(_03616_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09481_ (.I(_03614_),
    .Z(_03617_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09482_ (.A1(\as2650.ivec[0] ),
    .A2(_03617_),
    .ZN(_03618_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09483_ (.A1(_01830_),
    .A2(_03616_),
    .B(_03618_),
    .ZN(_00275_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09484_ (.A1(\as2650.ivec[1] ),
    .A2(_03617_),
    .ZN(_03619_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09485_ (.A1(_01851_),
    .A2(_03616_),
    .B(_03619_),
    .ZN(_00276_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09486_ (.I0(\as2650.ivec[2] ),
    .I1(_02067_),
    .S(_03615_),
    .Z(_03620_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09487_ (.I(_03620_),
    .Z(_00277_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09488_ (.I0(\as2650.ivec[3] ),
    .I1(_02098_),
    .S(_03615_),
    .Z(_03621_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09489_ (.I(_03621_),
    .Z(_00278_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09490_ (.I(_02120_),
    .Z(_03622_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09491_ (.I0(\as2650.ivec[4] ),
    .I1(_03622_),
    .S(_03615_),
    .Z(_03623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09492_ (.I(_03623_),
    .Z(_00279_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09493_ (.A1(\as2650.ivec[5] ),
    .A2(_03617_),
    .ZN(_03624_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09494_ (.A1(_01900_),
    .A2(_03616_),
    .B(_03624_),
    .ZN(_00280_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09495_ (.I(_01911_),
    .Z(_03625_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09496_ (.A1(\as2650.ivec[6] ),
    .A2(_03617_),
    .ZN(_03626_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09497_ (.A1(_03625_),
    .A2(_03616_),
    .B(_03626_),
    .ZN(_00281_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09498_ (.I0(\as2650.ivec[7] ),
    .I1(_03285_),
    .S(_03614_),
    .Z(_03627_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09499_ (.I(_03627_),
    .Z(_00282_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09500_ (.I(_02686_),
    .Z(_03628_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09501_ (.I(_03628_),
    .Z(_03629_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09502_ (.A1(_03510_),
    .A2(_02255_),
    .A3(_02402_),
    .ZN(_03630_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09503_ (.I(_03630_),
    .Z(_03631_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09504_ (.A1(\as2650.stack[2][0] ),
    .A2(_03631_),
    .ZN(_03632_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09505_ (.A1(_01840_),
    .A2(_02697_),
    .B(_02699_),
    .ZN(_03633_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09506_ (.A1(_03557_),
    .A2(_03629_),
    .B1(_03632_),
    .B2(_03633_),
    .ZN(_00283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09507_ (.A1(\as2650.stack[2][1] ),
    .A2(_03631_),
    .ZN(_03634_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09508_ (.I(_02681_),
    .Z(_03635_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09509_ (.I(_02687_),
    .Z(_03636_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09510_ (.A1(_01858_),
    .A2(_03635_),
    .B(_03636_),
    .ZN(_03637_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09511_ (.A1(_03564_),
    .A2(_03629_),
    .B1(_03634_),
    .B2(_03637_),
    .ZN(_00284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09512_ (.A1(\as2650.stack[2][2] ),
    .A2(_03631_),
    .ZN(_03638_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09513_ (.A1(_01870_),
    .A2(_03635_),
    .B(_03636_),
    .ZN(_03639_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09514_ (.A1(_03569_),
    .A2(_03629_),
    .B1(_03638_),
    .B2(_03639_),
    .ZN(_00285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09515_ (.A1(\as2650.stack[2][3] ),
    .A2(_03631_),
    .ZN(_03640_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09516_ (.A1(_01881_),
    .A2(_03635_),
    .B(_03636_),
    .ZN(_03641_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09517_ (.A1(_03572_),
    .A2(_03629_),
    .B1(_03640_),
    .B2(_03641_),
    .ZN(_00286_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09518_ (.I(_02687_),
    .Z(_03642_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09519_ (.I(_03630_),
    .Z(_03643_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09520_ (.A1(\as2650.stack[2][4] ),
    .A2(_03643_),
    .ZN(_03644_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09521_ (.A1(_01892_),
    .A2(_03635_),
    .B(_03636_),
    .ZN(_03645_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09522_ (.A1(_03575_),
    .A2(_03642_),
    .B1(_03644_),
    .B2(_03645_),
    .ZN(_00287_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09523_ (.A1(\as2650.stack[2][5] ),
    .A2(_03643_),
    .ZN(_03646_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09524_ (.A1(_01906_),
    .A2(_02684_),
    .B(_03628_),
    .ZN(_03647_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09525_ (.A1(_03580_),
    .A2(_03642_),
    .B1(_03646_),
    .B2(_03647_),
    .ZN(_00288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09526_ (.A1(\as2650.stack[2][6] ),
    .A2(_03643_),
    .ZN(_03648_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09527_ (.A1(_01916_),
    .A2(_02684_),
    .B(_03628_),
    .ZN(_03649_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09528_ (.A1(_03583_),
    .A2(_03642_),
    .B1(_03648_),
    .B2(_03649_),
    .ZN(_00289_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09529_ (.A1(\as2650.stack[2][7] ),
    .A2(_03643_),
    .ZN(_03650_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09530_ (.A1(_01925_),
    .A2(_02684_),
    .B(_03628_),
    .ZN(_03651_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09531_ (.A1(_03586_),
    .A2(_03642_),
    .B1(_03650_),
    .B2(_03651_),
    .ZN(_00290_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09532_ (.A1(_00705_),
    .A2(_00681_),
    .ZN(_03652_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09533_ (.A1(_00875_),
    .A2(_00825_),
    .ZN(_03653_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09534_ (.I(_02901_),
    .Z(_03654_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _09535_ (.A1(_00832_),
    .A2(_00905_),
    .ZN(_03655_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09536_ (.I(_03655_),
    .Z(_03656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _09537_ (.A1(_02747_),
    .A2(_03655_),
    .ZN(_03657_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09538_ (.A1(_00466_),
    .A2(_00907_),
    .A3(_02331_),
    .A4(_03657_),
    .ZN(_03658_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09539_ (.A1(_03654_),
    .A2(_03656_),
    .B(_03658_),
    .ZN(_03659_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09540_ (.A1(_00906_),
    .A2(_02334_),
    .B(_00894_),
    .ZN(_03660_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _09541_ (.A1(_03652_),
    .A2(_03653_),
    .B(_03659_),
    .C(_03660_),
    .ZN(_03661_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09542_ (.I(_02750_),
    .Z(_03662_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09543_ (.I(_03662_),
    .Z(_03663_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09544_ (.A1(_00642_),
    .A2(_00580_),
    .ZN(_03664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09545_ (.A1(_00928_),
    .A2(_03664_),
    .ZN(_03665_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09546_ (.I(_03653_),
    .Z(_03666_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _09547_ (.A1(_03663_),
    .A2(_03665_),
    .B(_03666_),
    .C(_00892_),
    .ZN(_03667_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09548_ (.A1(_00696_),
    .A2(_00532_),
    .A3(\as2650.cycle[4] ),
    .ZN(_03668_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09549_ (.A1(_00625_),
    .A2(_00647_),
    .ZN(_03669_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09550_ (.A1(_03668_),
    .A2(_03669_),
    .Z(_03670_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09551_ (.I(_03670_),
    .Z(_03671_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09552_ (.A1(_00804_),
    .A2(_01016_),
    .A3(\as2650.cycle[4] ),
    .ZN(_03672_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09553_ (.A1(_00679_),
    .A2(_00533_),
    .ZN(_03673_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09554_ (.A1(_01033_),
    .A2(_03673_),
    .ZN(_03674_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _09555_ (.I(_03674_),
    .ZN(_03675_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09556_ (.A1(_00709_),
    .A2(_03675_),
    .B(_00837_),
    .ZN(_03676_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09557_ (.A1(_00483_),
    .A2(_03672_),
    .B(_03676_),
    .ZN(_03677_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _09558_ (.A1(_03661_),
    .A2(_03667_),
    .A3(_03671_),
    .A4(_03677_),
    .ZN(_03678_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09559_ (.I(_00627_),
    .Z(_03679_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09560_ (.I(_03679_),
    .Z(_03680_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09561_ (.I(_00628_),
    .Z(_03681_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09562_ (.A1(_03681_),
    .A2(_00844_),
    .ZN(_03682_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09563_ (.A1(_03680_),
    .A2(_00713_),
    .B(_03682_),
    .ZN(_03683_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09564_ (.A1(net26),
    .A2(_03678_),
    .B(_00883_),
    .ZN(_03684_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09565_ (.A1(_03678_),
    .A2(_03683_),
    .B(_03684_),
    .ZN(_00291_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09566_ (.I(_02525_),
    .Z(_03685_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09567_ (.A1(_00954_),
    .A2(_00705_),
    .A3(_03685_),
    .ZN(_03686_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09568_ (.A1(net24),
    .A2(_03686_),
    .ZN(_03687_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09569_ (.I(_00909_),
    .Z(_03688_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09570_ (.I(_03688_),
    .Z(_03689_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09571_ (.A1(_01118_),
    .A2(_03686_),
    .B(_03687_),
    .C(_03689_),
    .ZN(_00292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09572_ (.A1(_00575_),
    .A2(_02508_),
    .ZN(_03690_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09573_ (.A1(_00642_),
    .A2(_02744_),
    .ZN(_03691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09574_ (.A1(_03664_),
    .A2(_02502_),
    .ZN(_03692_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09575_ (.I(_00698_),
    .Z(_03693_));
 gf180mcu_fd_sc_mcu7t5v0__oai33_1 _09576_ (.A1(_00502_),
    .A2(_03690_),
    .A3(_03691_),
    .B1(_03692_),
    .B2(_00725_),
    .B3(_03693_),
    .ZN(_03694_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09577_ (.I(net83),
    .ZN(_03695_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _09578_ (.A1(_00967_),
    .A2(_02519_),
    .B(_03695_),
    .C(_00692_),
    .ZN(_03696_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09579_ (.I(_03656_),
    .Z(_03697_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09580_ (.A1(_02903_),
    .A2(_00675_),
    .A3(_03697_),
    .ZN(_03698_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09581_ (.A1(_00497_),
    .A2(_00705_),
    .B(_02537_),
    .ZN(_03699_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09582_ (.A1(_03690_),
    .A2(_03698_),
    .B(_03699_),
    .ZN(_03700_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09583_ (.A1(_03696_),
    .A2(_03700_),
    .B(net25),
    .ZN(_03701_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09584_ (.I(_00506_),
    .Z(_03702_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09585_ (.I(_02486_),
    .Z(_03703_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _09586_ (.A1(_00576_),
    .A2(_03703_),
    .B(_03696_),
    .C(_03700_),
    .ZN(_03704_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09587_ (.A1(_03702_),
    .A2(_03704_),
    .ZN(_03705_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09588_ (.A1(_03701_),
    .A2(_03705_),
    .ZN(_00293_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _09589_ (.A1(_00459_),
    .A2(_00715_),
    .A3(_00518_),
    .A4(_03685_),
    .ZN(_03706_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09590_ (.A1(_00944_),
    .A2(_02487_),
    .ZN(_03707_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _09591_ (.A1(_00650_),
    .A2(_00822_),
    .A3(_03685_),
    .ZN(_03708_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09592_ (.A1(_02515_),
    .A2(_02519_),
    .ZN(_03709_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _09593_ (.A1(_00716_),
    .A2(_00855_),
    .A3(_03709_),
    .ZN(_03710_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _09594_ (.A1(_02565_),
    .A2(_02500_),
    .B(_03708_),
    .C(_03710_),
    .ZN(_03711_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09595_ (.A1(_00946_),
    .A2(_00948_),
    .A3(_00903_),
    .ZN(_03712_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09596_ (.A1(_02744_),
    .A2(_00978_),
    .ZN(_03713_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _09597_ (.A1(_00966_),
    .A2(_03712_),
    .A3(_03685_),
    .A4(_03713_),
    .ZN(_03714_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09598_ (.A1(_02526_),
    .A2(_03714_),
    .ZN(_03715_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09599_ (.A1(_00905_),
    .A2(_00822_),
    .A3(_02486_),
    .ZN(_03716_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _09600_ (.A1(_00828_),
    .A2(_00954_),
    .A3(_03716_),
    .ZN(_03717_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09601_ (.A1(_02533_),
    .A2(_02541_),
    .A3(_03717_),
    .ZN(_03718_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _09602_ (.A1(_03707_),
    .A2(_03711_),
    .A3(_03715_),
    .A4(_03718_),
    .ZN(_03719_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09603_ (.A1(_00798_),
    .A2(_00654_),
    .A3(_03668_),
    .ZN(_03720_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _09604_ (.A1(_00759_),
    .A2(_03720_),
    .ZN(_03721_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09605_ (.A1(_00634_),
    .A2(_00768_),
    .B(_00633_),
    .ZN(_03722_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09606_ (.A1(_03722_),
    .A2(_00637_),
    .ZN(_03723_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09607_ (.A1(_00607_),
    .A2(_03723_),
    .ZN(_03724_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _09608_ (.A1(_00781_),
    .A2(_00759_),
    .A3(_03672_),
    .Z(_03725_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09609_ (.A1(_02523_),
    .A2(_03725_),
    .ZN(_03726_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09610_ (.A1(_03721_),
    .A2(_03724_),
    .B(_03726_),
    .ZN(_03727_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09611_ (.I(_02508_),
    .Z(_03728_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09612_ (.I(_03728_),
    .Z(_03729_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09613_ (.A1(_00665_),
    .A2(_03729_),
    .ZN(_03730_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09614_ (.A1(_02535_),
    .A2(_02540_),
    .B(_02532_),
    .ZN(_03731_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09615_ (.A1(_00799_),
    .A2(_00623_),
    .A3(_01793_),
    .ZN(_03732_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _09616_ (.A1(net84),
    .A2(_00473_),
    .A3(_00546_),
    .A4(_03703_),
    .ZN(_03733_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _09617_ (.A1(_03730_),
    .A2(_03731_),
    .A3(_03732_),
    .A4(_03733_),
    .Z(_03734_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09618_ (.A1(_00758_),
    .A2(_00916_),
    .A3(_03728_),
    .ZN(_03735_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09619_ (.I(_01790_),
    .Z(_03736_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09620_ (.A1(_00912_),
    .A2(_00495_),
    .B(_02332_),
    .ZN(_03737_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _09621_ (.A1(_00691_),
    .A2(_03736_),
    .B(_03737_),
    .ZN(_03738_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _09622_ (.A1(_00799_),
    .A2(_00967_),
    .B1(_00760_),
    .B2(_03735_),
    .C(_03738_),
    .ZN(_03739_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09623_ (.A1(_00660_),
    .A2(_02508_),
    .ZN(_03740_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09624_ (.A1(_01791_),
    .A2(_02493_),
    .ZN(_03741_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _09625_ (.A1(_01033_),
    .A2(_00873_),
    .A3(_02514_),
    .A4(_02519_),
    .ZN(_03742_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09626_ (.A1(_00703_),
    .A2(_03740_),
    .B(_03741_),
    .C(_03742_),
    .ZN(_03743_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09627_ (.A1(_03739_),
    .A2(_03743_),
    .ZN(_03744_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _09628_ (.A1(_03727_),
    .A2(_03734_),
    .A3(_03744_),
    .ZN(_03745_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _09629_ (.A1(_02504_),
    .A2(_03706_),
    .A3(_03719_),
    .A4(_03745_),
    .ZN(_03746_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09630_ (.I(_03746_),
    .Z(_03747_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09631_ (.I(_03747_),
    .Z(_03748_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09632_ (.A1(_00825_),
    .A2(_02560_),
    .ZN(_03749_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _09633_ (.A1(_00969_),
    .A2(_03749_),
    .ZN(_03750_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09634_ (.I(_03750_),
    .Z(_03751_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _09635_ (.I(net55),
    .ZN(_03752_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09636_ (.I(_03752_),
    .Z(_03753_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09637_ (.I(_00833_),
    .Z(_03754_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09638_ (.I(_01705_),
    .Z(_03755_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09639_ (.I(_03755_),
    .Z(_03756_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09640_ (.I(_03756_),
    .Z(_03757_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _09641_ (.A1(_03752_),
    .A2(_03109_),
    .Z(_03758_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09642_ (.I(net100),
    .Z(_03759_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09643_ (.I(_03755_),
    .Z(_03760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09644_ (.A1(_03759_),
    .A2(_03760_),
    .ZN(_03761_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09645_ (.I(_00918_),
    .Z(_03762_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _09646_ (.A1(_00830_),
    .A2(_03762_),
    .A3(_00732_),
    .ZN(_03763_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09647_ (.A1(_03757_),
    .A2(_03758_),
    .B(_03761_),
    .C(_03763_),
    .ZN(_03764_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09648_ (.I(_01834_),
    .Z(_03765_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09649_ (.A1(_00828_),
    .A2(_00858_),
    .ZN(_03766_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09650_ (.A1(_03765_),
    .A2(_03766_),
    .ZN(_03767_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09651_ (.I(_03109_),
    .Z(_03768_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09652_ (.A1(_00629_),
    .A2(_03693_),
    .Z(_03769_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09653_ (.I(_03769_),
    .Z(_03770_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09654_ (.A1(_00629_),
    .A2(_00661_),
    .ZN(_03771_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09655_ (.I(_03771_),
    .Z(_03772_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09656_ (.I(_00699_),
    .Z(_03773_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09657_ (.A1(_03759_),
    .A2(_03773_),
    .B(_02515_),
    .ZN(_03774_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09658_ (.A1(_03768_),
    .A2(_03770_),
    .B1(_03772_),
    .B2(_03759_),
    .C(_03774_),
    .ZN(_03775_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09659_ (.A1(_03767_),
    .A2(_03775_),
    .B(_00718_),
    .ZN(_03776_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09660_ (.A1(_03752_),
    .A2(_02549_),
    .ZN(_03777_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _09661_ (.A1(_03754_),
    .A2(_03764_),
    .A3(_03776_),
    .A4(_03777_),
    .ZN(_03778_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09662_ (.A1(_03753_),
    .A2(_00834_),
    .B(_03679_),
    .C(_03778_),
    .ZN(_03779_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09663_ (.I(_00597_),
    .Z(_03780_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09664_ (.I(net100),
    .ZN(_03781_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09665_ (.A1(_00754_),
    .A2(_00770_),
    .ZN(_03782_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09666_ (.I(_03782_),
    .Z(_03783_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09667_ (.A1(_03089_),
    .A2(_01094_),
    .Z(_03784_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09668_ (.I(_00769_),
    .Z(_03785_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09669_ (.A1(_02856_),
    .A2(_03784_),
    .B(_03785_),
    .ZN(_03786_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09670_ (.A1(_03768_),
    .A2(_03784_),
    .B(_03786_),
    .ZN(_03787_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09671_ (.I(_01026_),
    .Z(_03788_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09672_ (.I(_03788_),
    .Z(_03789_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _09673_ (.A1(_01078_),
    .A2(_01050_),
    .ZN(_03790_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09674_ (.I(_01103_),
    .Z(_03791_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09675_ (.I(_03791_),
    .Z(_03792_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09676_ (.A1(_03792_),
    .A2(_01051_),
    .Z(_03793_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09677_ (.I(_03722_),
    .Z(_03794_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _09678_ (.A1(_03789_),
    .A2(_03790_),
    .B1(_03793_),
    .B2(_03768_),
    .C(_03794_),
    .ZN(_03795_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09679_ (.A1(_03787_),
    .A2(_03795_),
    .ZN(_03796_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09680_ (.I(_00755_),
    .Z(_03797_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09681_ (.A1(_03781_),
    .A2(_03783_),
    .B1(_03796_),
    .B2(_03797_),
    .ZN(_03798_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09682_ (.A1(_00598_),
    .A2(_03758_),
    .ZN(_03799_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09683_ (.I(_03673_),
    .Z(_03800_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09684_ (.I(_03800_),
    .Z(_03801_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09685_ (.A1(_03780_),
    .A2(_03798_),
    .B(_03799_),
    .C(_03801_),
    .ZN(_03802_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09686_ (.A1(_03779_),
    .A2(_03802_),
    .ZN(_03803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09687_ (.A1(_00777_),
    .A2(_03803_),
    .ZN(_03804_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09688_ (.A1(_01836_),
    .A2(_03751_),
    .B(_03804_),
    .ZN(_03805_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09689_ (.I(_03746_),
    .Z(_03806_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09690_ (.I(_03806_),
    .Z(_03807_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09691_ (.A1(_03759_),
    .A2(_03807_),
    .B(_00883_),
    .ZN(_03808_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09692_ (.A1(_03748_),
    .A2(_03805_),
    .B(_03808_),
    .ZN(_00294_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _09693_ (.I(_01853_),
    .ZN(_03809_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09694_ (.I(_03656_),
    .Z(_03810_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09695_ (.A1(_00526_),
    .A2(_00708_),
    .ZN(_03811_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09696_ (.I(_03811_),
    .Z(_03812_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09697_ (.A1(_00919_),
    .A2(_03812_),
    .ZN(_03813_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09698_ (.A1(_00829_),
    .A2(_00732_),
    .ZN(_03814_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09699_ (.I(_03814_),
    .Z(_03815_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09700_ (.I(net31),
    .Z(_03816_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09701_ (.I(_00848_),
    .Z(_03817_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09702_ (.I(_03817_),
    .Z(_03818_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09703_ (.A1(net55),
    .A2(net8),
    .ZN(_03819_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_4 _09704_ (.A1(net56),
    .A2(net9),
    .ZN(_03820_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09705_ (.A1(_03819_),
    .A2(_03820_),
    .ZN(_03821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09706_ (.A1(_00850_),
    .A2(_03821_),
    .ZN(_03822_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09707_ (.A1(_03816_),
    .A2(_03818_),
    .B(_03822_),
    .ZN(_03823_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09708_ (.I(_03769_),
    .Z(_03824_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09709_ (.I(_03771_),
    .Z(_03825_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09710_ (.I(_03825_),
    .Z(_03826_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09711_ (.I(_00723_),
    .Z(_03827_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _09712_ (.A1(net31),
    .A2(_03781_),
    .Z(_03828_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09713_ (.A1(_03827_),
    .A2(_03828_),
    .ZN(_03829_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09714_ (.A1(_02858_),
    .A2(_03824_),
    .B1(_03826_),
    .B2(_03816_),
    .C(_03829_),
    .ZN(_03830_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09715_ (.A1(_03815_),
    .A2(_03823_),
    .B1(_03830_),
    .B2(_00734_),
    .ZN(_03831_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09716_ (.I(_03762_),
    .Z(_03832_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09717_ (.I(_03832_),
    .Z(_03833_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09718_ (.A1(_01855_),
    .A2(_03813_),
    .B1(_03831_),
    .B2(_03833_),
    .ZN(_03834_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09719_ (.I(_00471_),
    .Z(_03835_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09720_ (.I(_03835_),
    .Z(_03836_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09721_ (.I(_03836_),
    .Z(_03837_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09722_ (.A1(_01834_),
    .A2(_01078_),
    .ZN(_03838_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09723_ (.A1(_03838_),
    .A2(_03820_),
    .Z(_03839_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09724_ (.I(_00635_),
    .Z(_03840_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _09725_ (.I(_01215_),
    .Z(_03841_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09726_ (.I(_01088_),
    .Z(_03842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09727_ (.A1(_01078_),
    .A2(_01093_),
    .ZN(_03843_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _09728_ (.A1(_05827_),
    .A2(_05833_),
    .ZN(_03844_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09729_ (.A1(_01213_),
    .A2(_03844_),
    .A3(_01203_),
    .Z(_03845_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09730_ (.A1(_03843_),
    .A2(_03845_),
    .ZN(_03846_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09731_ (.A1(_03843_),
    .A2(_03845_),
    .ZN(_03847_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09732_ (.A1(_03842_),
    .A2(_03847_),
    .ZN(_03848_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09733_ (.A1(_03841_),
    .A2(_03842_),
    .B1(_03846_),
    .B2(_03848_),
    .ZN(_03849_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _09734_ (.A1(_01213_),
    .A2(_03844_),
    .A3(_01196_),
    .Z(_03850_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09735_ (.A1(_03790_),
    .A2(_03850_),
    .B(_03791_),
    .ZN(_03851_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09736_ (.A1(_03790_),
    .A2(_03850_),
    .B(_03851_),
    .ZN(_03852_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09737_ (.A1(_03841_),
    .A2(_03788_),
    .B(_03852_),
    .ZN(_03853_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09738_ (.A1(_03840_),
    .A2(_03849_),
    .B1(_03853_),
    .B2(_03794_),
    .ZN(_03854_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09739_ (.A1(_00618_),
    .A2(_03854_),
    .ZN(_03855_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _09740_ (.A1(_03782_),
    .A2(_03828_),
    .B(_03855_),
    .C(_00865_),
    .ZN(_03856_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09741_ (.I(_00906_),
    .Z(_03857_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09742_ (.I(_02559_),
    .Z(_03858_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09743_ (.A1(_03857_),
    .A2(_03858_),
    .ZN(_03859_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _09744_ (.A1(_03780_),
    .A2(_03839_),
    .B(_03856_),
    .C(_03859_),
    .ZN(_03860_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09745_ (.A1(_03809_),
    .A2(_03810_),
    .B1(_03834_),
    .B2(_03837_),
    .C(_03860_),
    .ZN(_03861_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _09746_ (.A1(_01855_),
    .A2(_03751_),
    .B1(_03861_),
    .B2(_02548_),
    .ZN(_03862_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09747_ (.I(_00845_),
    .Z(_03863_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09748_ (.A1(_03816_),
    .A2(_03807_),
    .B(_03863_),
    .ZN(_03864_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09749_ (.A1(_03748_),
    .A2(_03862_),
    .B(_03864_),
    .ZN(_00295_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09750_ (.I(_00775_),
    .Z(_03865_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09751_ (.I(_00907_),
    .Z(_03866_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09752_ (.A1(_03865_),
    .A2(_03866_),
    .ZN(_03867_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09753_ (.I(_03859_),
    .Z(_03868_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _09754_ (.A1(net57),
    .A2(net10),
    .ZN(_03869_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _09755_ (.A1(net56),
    .A2(_01214_),
    .ZN(_03870_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09756_ (.A1(_03838_),
    .A2(_03820_),
    .B(_03870_),
    .ZN(_03871_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09757_ (.A1(_03869_),
    .A2(_03871_),
    .Z(_03872_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09758_ (.I(_03782_),
    .Z(_03873_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09759_ (.I(net99),
    .ZN(_03874_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09760_ (.A1(_03816_),
    .A2(net100),
    .ZN(_03875_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09761_ (.A1(_03874_),
    .A2(_03875_),
    .Z(_03876_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09762_ (.I(_03089_),
    .Z(_03877_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09763_ (.A1(_01216_),
    .A2(_01206_),
    .B(_03847_),
    .ZN(_03878_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09764_ (.A1(_01264_),
    .A2(_01260_),
    .Z(_03879_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09765_ (.A1(_03878_),
    .A2(_03879_),
    .B(_03842_),
    .ZN(_03880_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09766_ (.A1(_03878_),
    .A2(_03879_),
    .B(_03880_),
    .ZN(_03881_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09767_ (.A1(_02860_),
    .A2(_03877_),
    .B(_03881_),
    .C(_03840_),
    .ZN(_03882_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09768_ (.I(_03788_),
    .Z(_03883_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09769_ (.I(_02925_),
    .Z(_03884_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09770_ (.I(_01213_),
    .ZN(_03885_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09771_ (.I(_03885_),
    .Z(_03886_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _09772_ (.A1(_03886_),
    .A2(_01197_),
    .A3(_01198_),
    .B1(_03790_),
    .B2(_03850_),
    .ZN(_03887_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09773_ (.A1(_03884_),
    .A2(_01254_),
    .A3(_03887_),
    .Z(_03888_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09774_ (.A1(_03884_),
    .A2(_03788_),
    .B(_00616_),
    .ZN(_03889_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09775_ (.A1(_03883_),
    .A2(_03888_),
    .B(_03889_),
    .ZN(_03890_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09776_ (.A1(_03882_),
    .A2(_03890_),
    .ZN(_03891_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09777_ (.I(_00755_),
    .Z(_03892_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09778_ (.A1(_03873_),
    .A2(_03876_),
    .B1(_03891_),
    .B2(_03892_),
    .ZN(_03893_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _09779_ (.I0(_03872_),
    .I1(_03893_),
    .S(_00610_),
    .Z(_03894_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09780_ (.A1(_00833_),
    .A2(_03813_),
    .ZN(_03895_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09781_ (.A1(_00716_),
    .A2(_00708_),
    .ZN(_03896_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09782_ (.I(_03773_),
    .Z(_03897_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09783_ (.I(_00786_),
    .Z(_03898_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09784_ (.I(_03898_),
    .Z(_03899_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09785_ (.A1(_02859_),
    .A2(_03899_),
    .ZN(_03900_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09786_ (.A1(_03874_),
    .A2(_00631_),
    .B1(_03772_),
    .B2(_03900_),
    .ZN(_03901_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09787_ (.A1(_03897_),
    .A2(_03876_),
    .B(_03901_),
    .C(_02561_),
    .ZN(_03902_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09788_ (.I(_02941_),
    .Z(_03903_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09789_ (.I(_00848_),
    .Z(_03904_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09790_ (.I(_03904_),
    .Z(_03905_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09791_ (.A1(_03819_),
    .A2(_03820_),
    .B(_03870_),
    .ZN(_03906_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09792_ (.A1(_03869_),
    .A2(_03906_),
    .Z(_03907_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09793_ (.A1(_03905_),
    .A2(_03907_),
    .ZN(_03908_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09794_ (.A1(net99),
    .A2(_03903_),
    .B(_03763_),
    .C(_03908_),
    .ZN(_03909_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09795_ (.A1(_03896_),
    .A2(_03902_),
    .B(_03909_),
    .ZN(_03910_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09796_ (.I(_00833_),
    .Z(_03911_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09797_ (.I(_03911_),
    .Z(_03912_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09798_ (.A1(_01868_),
    .A2(_03895_),
    .B1(_03910_),
    .B2(_03912_),
    .ZN(_03913_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09799_ (.I(_00906_),
    .Z(_03914_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09800_ (.I(_03914_),
    .Z(_03915_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09801_ (.A1(_03868_),
    .A2(_03894_),
    .B1(_03913_),
    .B2(_03915_),
    .ZN(_03916_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09802_ (.I(_00776_),
    .Z(_03917_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09803_ (.A1(_01868_),
    .A2(_03867_),
    .B1(_03916_),
    .B2(_03917_),
    .ZN(_03918_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09804_ (.A1(net99),
    .A2(_03807_),
    .B(_03863_),
    .ZN(_03919_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09805_ (.A1(_03748_),
    .A2(_03918_),
    .B(_03919_),
    .ZN(_00296_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09806_ (.I(net58),
    .Z(_03920_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09807_ (.I(_03920_),
    .Z(_03921_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09808_ (.I(_03750_),
    .Z(_03922_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09809_ (.I(_00875_),
    .Z(_03923_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09810_ (.I(_03811_),
    .Z(_03924_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09811_ (.I(_03924_),
    .Z(_03925_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _09812_ (.A1(_03923_),
    .A2(_00794_),
    .A3(_03925_),
    .ZN(_03926_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09813_ (.I(_03858_),
    .Z(_03927_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09814_ (.A1(_03911_),
    .A2(_03927_),
    .ZN(_03928_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09815_ (.A1(_03920_),
    .A2(_02861_),
    .ZN(_03929_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09816_ (.I(_03929_),
    .ZN(_03930_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09817_ (.A1(_03920_),
    .A2(_02861_),
    .ZN(_03931_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09818_ (.A1(_03930_),
    .A2(_03931_),
    .ZN(_03932_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09819_ (.A1(_01866_),
    .A2(_01264_),
    .ZN(_03933_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09820_ (.I(_03869_),
    .ZN(_03934_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09821_ (.A1(_03934_),
    .A2(_03906_),
    .ZN(_03935_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09822_ (.A1(_03933_),
    .A2(_03935_),
    .Z(_03936_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09823_ (.A1(_03932_),
    .A2(_03936_),
    .ZN(_03937_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09824_ (.A1(_03905_),
    .A2(_03937_),
    .ZN(_03938_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09825_ (.A1(net98),
    .A2(_00604_),
    .B(_03938_),
    .ZN(_03939_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _09826_ (.I(net98),
    .ZN(_03940_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _09827_ (.A1(net99),
    .A2(net31),
    .A3(net100),
    .ZN(_03941_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09828_ (.A1(_03940_),
    .A2(_03941_),
    .Z(_03942_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09829_ (.A1(_00928_),
    .A2(_03942_),
    .ZN(_03943_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _09830_ (.A1(_02864_),
    .A2(_03824_),
    .B1(_03826_),
    .B2(net98),
    .C(_03896_),
    .ZN(_03944_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09831_ (.A1(_03815_),
    .A2(_03939_),
    .B1(_03943_),
    .B2(_03944_),
    .ZN(_03945_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09832_ (.A1(_03921_),
    .A2(_03926_),
    .B1(_03928_),
    .B2(_03945_),
    .ZN(_03946_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09833_ (.I(_00865_),
    .Z(_03947_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09834_ (.A1(_03934_),
    .A2(_03871_),
    .ZN(_03948_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09835_ (.A1(_03933_),
    .A2(_03948_),
    .Z(_03949_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09836_ (.A1(_03932_),
    .A2(_03949_),
    .Z(_03950_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09837_ (.I(_01328_),
    .Z(_03951_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _09838_ (.A1(_03886_),
    .A2(_01204_),
    .A3(_01205_),
    .B1(_03843_),
    .B2(_03845_),
    .ZN(_03952_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09839_ (.A1(_01255_),
    .A2(_01259_),
    .B(_02924_),
    .ZN(_03953_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _09840_ (.A1(_02924_),
    .A2(_01255_),
    .A3(_01259_),
    .ZN(_03954_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09841_ (.A1(_03952_),
    .A2(_03953_),
    .B(_03954_),
    .ZN(_03955_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09842_ (.A1(_01528_),
    .A2(_01320_),
    .ZN(_03956_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09843_ (.A1(_01262_),
    .A2(_01527_),
    .B1(_01321_),
    .B2(_01322_),
    .ZN(_03957_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09844_ (.A1(_03956_),
    .A2(_03957_),
    .ZN(_03958_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09845_ (.A1(_01328_),
    .A2(_03958_),
    .ZN(_03959_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09846_ (.I(_02861_),
    .Z(_03960_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09847_ (.A1(_03960_),
    .A2(_01323_),
    .ZN(_03961_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09848_ (.A1(_03959_),
    .A2(_03961_),
    .ZN(_03962_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09849_ (.A1(_03955_),
    .A2(_03962_),
    .B(_03842_),
    .ZN(_03963_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09850_ (.A1(_03955_),
    .A2(_03962_),
    .B(_03963_),
    .ZN(_03964_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09851_ (.A1(_03951_),
    .A2(_03877_),
    .B(_03964_),
    .C(_00636_),
    .ZN(_03965_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09852_ (.A1(_01243_),
    .A2(_01248_),
    .B(_01253_),
    .C(_02925_),
    .ZN(_03966_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09853_ (.A1(_01251_),
    .A2(_01252_),
    .B(_01405_),
    .ZN(_03967_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _09854_ (.A1(_01405_),
    .A2(_01248_),
    .B(_03967_),
    .C(_02925_),
    .ZN(_03968_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09855_ (.A1(_03887_),
    .A2(_03966_),
    .B(_03968_),
    .ZN(_03969_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _09856_ (.A1(_02863_),
    .A2(_01343_),
    .A3(_03969_),
    .Z(_03970_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09857_ (.A1(_02864_),
    .A2(_03789_),
    .ZN(_03971_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09858_ (.I(_03794_),
    .Z(_03972_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _09859_ (.A1(_03883_),
    .A2(_03970_),
    .B(_03971_),
    .C(_03972_),
    .ZN(_03973_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09860_ (.A1(_03965_),
    .A2(_03973_),
    .B(_00766_),
    .ZN(_03974_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09861_ (.A1(_00755_),
    .A2(_00770_),
    .Z(_03975_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09862_ (.A1(_03975_),
    .A2(_03942_),
    .B(_00610_),
    .ZN(_03976_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09863_ (.A1(_03974_),
    .A2(_03976_),
    .ZN(_03977_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09864_ (.A1(_03947_),
    .A2(_03950_),
    .B(_03977_),
    .ZN(_03978_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09865_ (.I(_03800_),
    .Z(_03979_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09866_ (.A1(_03681_),
    .A2(_03946_),
    .B1(_03978_),
    .B2(_03979_),
    .ZN(_03980_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09867_ (.I(_00969_),
    .Z(_03981_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09868_ (.I(_03981_),
    .Z(_03982_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09869_ (.A1(_03921_),
    .A2(_03922_),
    .B1(_03980_),
    .B2(_03982_),
    .ZN(_03983_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09870_ (.I(_03806_),
    .Z(_03984_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09871_ (.A1(net98),
    .A2(_03984_),
    .B(_03863_),
    .ZN(_03985_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09872_ (.A1(_03748_),
    .A2(_03983_),
    .B(_03985_),
    .ZN(_00297_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09873_ (.I(_03702_),
    .Z(_03986_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09874_ (.I(_03750_),
    .Z(_03987_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09875_ (.I(net60),
    .Z(_03988_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09876_ (.A1(_03988_),
    .A2(net12),
    .Z(_03989_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _09877_ (.I(_03989_),
    .Z(_03990_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09878_ (.A1(_03929_),
    .A2(_03949_),
    .B(_03931_),
    .ZN(_03991_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09879_ (.A1(_03990_),
    .A2(_03991_),
    .Z(_03992_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09880_ (.A1(_03990_),
    .A2(_03991_),
    .B(_00597_),
    .ZN(_03993_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09881_ (.A1(_03940_),
    .A2(_03941_),
    .ZN(_03994_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09882_ (.A1(net97),
    .A2(_03994_),
    .Z(_03995_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09883_ (.A1(_01423_),
    .A2(_01412_),
    .Z(_03996_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09884_ (.A1(_01341_),
    .A2(_01342_),
    .B(_03960_),
    .ZN(_03997_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _09885_ (.A1(_03960_),
    .A2(_01341_),
    .A3(_01342_),
    .ZN(_03998_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09886_ (.A1(_03969_),
    .A2(_03997_),
    .B(_03998_),
    .ZN(_03999_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09887_ (.A1(_03996_),
    .A2(_03999_),
    .Z(_04000_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09888_ (.A1(_03996_),
    .A2(_03999_),
    .B(_03791_),
    .ZN(_04001_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _09889_ (.A1(_02915_),
    .A2(_03792_),
    .B1(_04000_),
    .B2(_04001_),
    .ZN(_04002_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09890_ (.I(_02915_),
    .Z(_04003_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09891_ (.A1(_01423_),
    .A2(_01415_),
    .Z(_04004_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09892_ (.A1(_03960_),
    .A2(_01323_),
    .ZN(_04005_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09893_ (.A1(_03955_),
    .A2(_04005_),
    .B(_03961_),
    .ZN(_04006_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09894_ (.A1(_04004_),
    .A2(_04006_),
    .B(_01088_),
    .ZN(_04007_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09895_ (.A1(_04004_),
    .A2(_04006_),
    .B(_04007_),
    .ZN(_04008_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09896_ (.A1(_04003_),
    .A2(_03089_),
    .B(_04008_),
    .ZN(_04009_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _09897_ (.A1(_03794_),
    .A2(_04002_),
    .B1(_04009_),
    .B2(_00635_),
    .ZN(_04010_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09898_ (.A1(_00618_),
    .A2(_04010_),
    .ZN(_04011_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09899_ (.A1(_03782_),
    .A2(_03995_),
    .B(_04011_),
    .ZN(_04012_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09900_ (.A1(_03992_),
    .A2(_03993_),
    .B1(_04012_),
    .B2(_00598_),
    .ZN(_04013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09901_ (.I(_03988_),
    .Z(_04014_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09902_ (.I(_04014_),
    .Z(_04015_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _09903_ (.A1(_00874_),
    .A2(_00532_),
    .ZN(_04016_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09904_ (.I(_04016_),
    .Z(_04017_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _09905_ (.I(net97),
    .ZN(_04018_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09906_ (.I(_00630_),
    .Z(_04019_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09907_ (.I(_03693_),
    .Z(_04020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09908_ (.A1(_00630_),
    .A2(_01426_),
    .ZN(_04021_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09909_ (.A1(_04018_),
    .A2(_04019_),
    .B(_04020_),
    .C(_04021_),
    .ZN(_04022_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09910_ (.A1(_00724_),
    .A2(_03995_),
    .B(_04022_),
    .C(_00733_),
    .ZN(_04023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09911_ (.I(_02932_),
    .Z(_04024_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09912_ (.A1(_03929_),
    .A2(_03936_),
    .B(_03931_),
    .ZN(_04025_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _09913_ (.A1(_03990_),
    .A2(_04025_),
    .ZN(_04026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09914_ (.A1(_04024_),
    .A2(_04026_),
    .ZN(_04027_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09915_ (.A1(net97),
    .A2(_00850_),
    .B(_03814_),
    .C(_04027_),
    .ZN(_04028_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09916_ (.A1(_04023_),
    .A2(_04028_),
    .ZN(_04029_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09917_ (.A1(_04015_),
    .A2(_03895_),
    .B1(_04017_),
    .B2(_04029_),
    .ZN(_04030_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09918_ (.I(_04030_),
    .ZN(_04031_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09919_ (.A1(_03801_),
    .A2(_04013_),
    .B1(_04031_),
    .B2(_03679_),
    .ZN(_04032_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09920_ (.I(_02547_),
    .Z(_04033_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _09921_ (.A1(_01889_),
    .A2(_03987_),
    .B1(_04032_),
    .B2(_04033_),
    .C(_03806_),
    .ZN(_04034_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09922_ (.A1(net97),
    .A2(_03807_),
    .B(_04034_),
    .ZN(_04035_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09923_ (.A1(_03986_),
    .A2(_04035_),
    .ZN(_00298_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09924_ (.I(_03747_),
    .Z(_04036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09925_ (.I(net35),
    .Z(_04037_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09926_ (.I(_03755_),
    .Z(_04038_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09927_ (.A1(net61),
    .A2(_02551_),
    .Z(_04039_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09928_ (.A1(_03990_),
    .A2(_04025_),
    .Z(_04040_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09929_ (.A1(_04014_),
    .A2(_01425_),
    .B(_04040_),
    .ZN(_04041_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09930_ (.A1(_04039_),
    .A2(_04041_),
    .Z(_04042_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09931_ (.A1(_03760_),
    .A2(_04042_),
    .ZN(_04043_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09932_ (.A1(_04037_),
    .A2(_04038_),
    .B(_04043_),
    .ZN(_04044_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _09933_ (.I(_02553_),
    .Z(_04045_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _09934_ (.A1(_04018_),
    .A2(_03940_),
    .A3(_03941_),
    .ZN(_04046_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09935_ (.A1(net35),
    .A2(_04046_),
    .Z(_04047_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09936_ (.I(_00661_),
    .Z(_04048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09937_ (.I(_04048_),
    .Z(_04049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _09938_ (.A1(_04045_),
    .A2(_03824_),
    .B1(_04047_),
    .B2(_04049_),
    .C1(_03826_),
    .C2(_04037_),
    .ZN(_04050_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09939_ (.A1(_03815_),
    .A2(_04044_),
    .B1(_04050_),
    .B2(_00734_),
    .ZN(_04051_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09940_ (.A1(_01903_),
    .A2(_03926_),
    .B1(_03928_),
    .B2(_04051_),
    .ZN(_04052_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09941_ (.A1(_01424_),
    .A2(_01413_),
    .Z(_04053_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09942_ (.A1(_03996_),
    .A2(_03999_),
    .B(_04053_),
    .ZN(_04054_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09943_ (.A1(_03203_),
    .A2(_01526_),
    .A3(_04054_),
    .Z(_04055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _09944_ (.A1(_03792_),
    .A2(_04055_),
    .ZN(_04056_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09945_ (.A1(_04045_),
    .A2(_03883_),
    .B(_00616_),
    .ZN(_04057_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09946_ (.A1(_01424_),
    .A2(_01416_),
    .Z(_04058_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09947_ (.A1(_04004_),
    .A2(_04006_),
    .B(_04058_),
    .ZN(_04059_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _09948_ (.A1(_01536_),
    .A2(_01531_),
    .A3(_04059_),
    .Z(_04060_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09949_ (.A1(_03877_),
    .A2(_04060_),
    .ZN(_04061_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09950_ (.I(_01088_),
    .Z(_04062_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09951_ (.I(_03785_),
    .Z(_04063_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09952_ (.A1(_04045_),
    .A2(_04062_),
    .B(_04063_),
    .ZN(_04064_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _09953_ (.A1(_04056_),
    .A2(_04057_),
    .B1(_04061_),
    .B2(_04064_),
    .ZN(_04065_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _09954_ (.A1(_03975_),
    .A2(_04047_),
    .B1(_04065_),
    .B2(_00766_),
    .C(_00764_),
    .ZN(_04066_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09955_ (.I(_04039_),
    .ZN(_04067_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09956_ (.A1(_04015_),
    .A2(_02849_),
    .B(_03992_),
    .ZN(_04068_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09957_ (.A1(_04067_),
    .A2(_04068_),
    .Z(_04069_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09958_ (.I(_03859_),
    .Z(_04070_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09959_ (.A1(_03947_),
    .A2(_04069_),
    .B(_04070_),
    .ZN(_04071_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09960_ (.A1(_03681_),
    .A2(_04052_),
    .B1(_04066_),
    .B2(_04071_),
    .ZN(_04072_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _09961_ (.A1(_01903_),
    .A2(_03922_),
    .B1(_04072_),
    .B2(_03982_),
    .ZN(_04073_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09962_ (.A1(_04037_),
    .A2(_03984_),
    .B(_03863_),
    .ZN(_04074_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09963_ (.A1(_04036_),
    .A2(_04073_),
    .B(_04074_),
    .ZN(_00299_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09964_ (.I(_04016_),
    .Z(_04075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _09965_ (.I(_03899_),
    .Z(_04076_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _09966_ (.I(net36),
    .Z(_04077_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09967_ (.A1(_04037_),
    .A2(_04046_),
    .ZN(_04078_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09968_ (.A1(_04077_),
    .A2(_04078_),
    .Z(_04079_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09969_ (.A1(_04076_),
    .A2(_04079_),
    .Z(_04080_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _09970_ (.A1(_02853_),
    .A2(_00721_),
    .B1(_00889_),
    .B2(_04077_),
    .C(_00733_),
    .ZN(_04081_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _09971_ (.I(_03817_),
    .Z(_04082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09972_ (.A1(net62),
    .A2(_01620_),
    .ZN(_04083_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _09973_ (.I(_04083_),
    .ZN(_04084_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09974_ (.A1(_01912_),
    .A2(_01620_),
    .ZN(_04085_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _09975_ (.A1(_04084_),
    .A2(_04085_),
    .ZN(_04086_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _09976_ (.I(net61),
    .ZN(_04087_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _09977_ (.A1(_03988_),
    .A2(net12),
    .B1(net1),
    .B2(_01901_),
    .ZN(_04088_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09978_ (.A1(_04087_),
    .A2(_01535_),
    .B(_04088_),
    .ZN(_04089_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _09979_ (.A1(_04040_),
    .A2(_04039_),
    .B(_04089_),
    .ZN(_04090_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _09980_ (.A1(_04086_),
    .A2(_04090_),
    .Z(_04091_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09981_ (.A1(_04082_),
    .A2(_04091_),
    .ZN(_04092_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _09982_ (.A1(_04077_),
    .A2(_02942_),
    .B(_03814_),
    .C(_04092_),
    .ZN(_04093_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09983_ (.A1(_04080_),
    .A2(_04081_),
    .B(_04093_),
    .ZN(_04094_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _09984_ (.A1(_01913_),
    .A2(_03895_),
    .B1(_04075_),
    .B2(_04094_),
    .C(_03915_),
    .ZN(_04095_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09985_ (.I(_01620_),
    .Z(_04096_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _09986_ (.A1(_04096_),
    .A2(_01630_),
    .Z(_04097_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09987_ (.A1(_02551_),
    .A2(_01530_),
    .ZN(_04098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09988_ (.A1(_02551_),
    .A2(_01530_),
    .ZN(_04099_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _09989_ (.A1(_04059_),
    .A2(_04098_),
    .B(_04099_),
    .ZN(_04100_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09990_ (.A1(_04097_),
    .A2(_04100_),
    .B(_03877_),
    .ZN(_04101_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _09991_ (.A1(_04097_),
    .A2(_04100_),
    .B(_04101_),
    .ZN(_04102_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _09992_ (.I(_03785_),
    .Z(_04103_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _09993_ (.A1(_02853_),
    .A2(_04062_),
    .B(_04102_),
    .C(_04103_),
    .ZN(_04104_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _09994_ (.A1(_01622_),
    .A2(_01613_),
    .Z(_04105_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _09995_ (.A1(_02552_),
    .A2(_01525_),
    .ZN(_04106_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _09996_ (.A1(_02552_),
    .A2(_01525_),
    .ZN(_04107_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _09997_ (.A1(_04054_),
    .A2(_04106_),
    .B(_04107_),
    .ZN(_04108_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _09998_ (.A1(_04105_),
    .A2(_04108_),
    .Z(_04109_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _09999_ (.A1(_04105_),
    .A2(_04108_),
    .B(_03792_),
    .ZN(_04110_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10000_ (.A1(_04109_),
    .A2(_04110_),
    .ZN(_04111_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10001_ (.I(_00616_),
    .Z(_04112_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _10002_ (.A1(_02854_),
    .A2(_03883_),
    .B(_04111_),
    .C(_04112_),
    .ZN(_04113_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _10003_ (.A1(_04104_),
    .A2(_04113_),
    .B(_03797_),
    .ZN(_04114_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10004_ (.A1(_03783_),
    .A2(_04079_),
    .B(_00598_),
    .ZN(_04115_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10005_ (.A1(_03992_),
    .A2(_04039_),
    .Z(_04116_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10006_ (.A1(_04089_),
    .A2(_04116_),
    .ZN(_04117_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10007_ (.A1(_04086_),
    .A2(_04117_),
    .ZN(_04118_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10008_ (.A1(_04114_),
    .A2(_04115_),
    .B1(_04118_),
    .B2(_00866_),
    .C(_04070_),
    .ZN(_04119_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10009_ (.A1(_04095_),
    .A2(_04119_),
    .B(_03865_),
    .ZN(_04120_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10010_ (.A1(_01913_),
    .A2(_03751_),
    .B(_04120_),
    .ZN(_04121_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10011_ (.I(_00845_),
    .Z(_04122_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10012_ (.A1(_04077_),
    .A2(_03984_),
    .B(_04122_),
    .ZN(_04123_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10013_ (.A1(_04036_),
    .A2(_04121_),
    .B(_04123_),
    .ZN(_00300_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10014_ (.I(_00826_),
    .Z(_04124_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10015_ (.I(_00718_),
    .Z(_04125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10016_ (.I(_03766_),
    .Z(_04126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10017_ (.I(net37),
    .Z(_04127_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10018_ (.A1(net36),
    .A2(net35),
    .A3(_04046_),
    .ZN(_04128_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10019_ (.A1(_04127_),
    .A2(_04128_),
    .Z(_04129_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10020_ (.A1(_03817_),
    .A2(_03770_),
    .B1(_03825_),
    .B2(_04127_),
    .C(_02748_),
    .ZN(_04130_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10021_ (.A1(_00724_),
    .A2(_04129_),
    .B(_04130_),
    .ZN(_04131_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10022_ (.A1(_01922_),
    .A2(_04126_),
    .B(_04131_),
    .ZN(_04132_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _10023_ (.I(net93),
    .ZN(_04133_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10024_ (.A1(_04133_),
    .A2(net2),
    .Z(_04134_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _10025_ (.I(_04134_),
    .ZN(_04135_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10026_ (.A1(_04085_),
    .A2(_04090_),
    .B(_04083_),
    .ZN(_04136_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10027_ (.A1(_04135_),
    .A2(_04136_),
    .Z(_04137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10028_ (.A1(_03903_),
    .A2(_04137_),
    .ZN(_04138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10029_ (.A1(_02560_),
    .A2(_03814_),
    .ZN(_04139_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10030_ (.A1(_04127_),
    .A2(_04038_),
    .B(_04139_),
    .ZN(_04140_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10031_ (.A1(_04125_),
    .A2(_04132_),
    .B1(_04138_),
    .B2(_04140_),
    .ZN(_04141_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10032_ (.I(_00876_),
    .Z(_04142_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10033_ (.A1(_01922_),
    .A2(_04017_),
    .B1(_04141_),
    .B2(_04142_),
    .ZN(_04143_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10034_ (.A1(_04085_),
    .A2(_04117_),
    .B(_04083_),
    .ZN(_04144_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10035_ (.A1(_04135_),
    .A2(_04144_),
    .Z(_04145_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _10036_ (.I(_04096_),
    .Z(_04146_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10037_ (.A1(_04146_),
    .A2(_01631_),
    .Z(_04147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10038_ (.A1(_04097_),
    .A2(_04100_),
    .B(_04147_),
    .ZN(_04148_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10039_ (.A1(_00601_),
    .A2(_01713_),
    .A3(_04148_),
    .Z(_04149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10040_ (.A1(_00603_),
    .A2(_04062_),
    .ZN(_04150_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10041_ (.A1(_04062_),
    .A2(_04149_),
    .B(_04150_),
    .C(_03840_),
    .ZN(_04151_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10042_ (.A1(_04146_),
    .A2(_01614_),
    .Z(_04152_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10043_ (.A1(_04152_),
    .A2(_04109_),
    .ZN(_04153_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _10044_ (.A1(_00601_),
    .A2(_01702_),
    .A3(_04153_),
    .Z(_04154_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10045_ (.A1(_00603_),
    .A2(_03789_),
    .ZN(_04155_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10046_ (.A1(_03789_),
    .A2(_04154_),
    .B(_04155_),
    .C(_03972_),
    .ZN(_04156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10047_ (.A1(_04151_),
    .A2(_04156_),
    .ZN(_04157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10048_ (.I(_00596_),
    .Z(_04158_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10049_ (.A1(_03783_),
    .A2(_04129_),
    .B1(_04157_),
    .B2(_03892_),
    .C(_04158_),
    .ZN(_04159_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10050_ (.A1(_03947_),
    .A2(_04145_),
    .B(_04159_),
    .ZN(_04160_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10051_ (.I(_03800_),
    .Z(_04161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10052_ (.A1(_04124_),
    .A2(_04143_),
    .B1(_04160_),
    .B2(_04161_),
    .ZN(_04162_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10053_ (.A1(_01922_),
    .A2(_03922_),
    .B1(_04162_),
    .B2(_03982_),
    .ZN(_04163_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10054_ (.A1(_04127_),
    .A2(_03984_),
    .B(_04122_),
    .ZN(_04164_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10055_ (.A1(_04036_),
    .A2(_04163_),
    .B(_04164_),
    .ZN(_00301_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10056_ (.I(net38),
    .Z(_04165_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10057_ (.A1(net64),
    .A2(_04096_),
    .Z(_04166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10058_ (.A1(_03989_),
    .A2(_04025_),
    .ZN(_04167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10059_ (.A1(_04086_),
    .A2(_04135_),
    .ZN(_04168_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10060_ (.I(_04168_),
    .ZN(_04169_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10061_ (.A1(net93),
    .A2(_01621_),
    .B1(_04089_),
    .B2(_04169_),
    .C(_04084_),
    .ZN(_04170_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _10062_ (.A1(_04167_),
    .A2(_04067_),
    .A3(_04168_),
    .B(_04170_),
    .ZN(_04171_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10063_ (.A1(_04166_),
    .A2(_04171_),
    .ZN(_04172_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10064_ (.A1(_03818_),
    .A2(_04172_),
    .ZN(_04173_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10065_ (.A1(_04165_),
    .A2(_02942_),
    .B(_03815_),
    .C(_04173_),
    .ZN(_04174_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10066_ (.I(net37),
    .ZN(_04175_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10067_ (.A1(_04175_),
    .A2(_04128_),
    .ZN(_04176_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10068_ (.A1(_04165_),
    .A2(_04176_),
    .Z(_04177_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10069_ (.I(_04165_),
    .ZN(_04178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10070_ (.I(\as2650.addr_buff[0] ),
    .Z(_04179_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10071_ (.A1(_04179_),
    .A2(_04048_),
    .ZN(_04180_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10072_ (.A1(_04178_),
    .A2(_00631_),
    .B1(_03772_),
    .B2(_04180_),
    .ZN(_04181_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10073_ (.A1(_00743_),
    .A2(_04177_),
    .B(_04181_),
    .C(_00734_),
    .ZN(_04182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10074_ (.A1(_04174_),
    .A2(_04182_),
    .ZN(_04183_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10075_ (.A1(_02185_),
    .A2(_03895_),
    .B1(_04017_),
    .B2(_04183_),
    .ZN(_04184_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10076_ (.I(\as2650.addr_buff[0] ),
    .ZN(_04185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10077_ (.I(_04185_),
    .Z(_04186_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _10078_ (.A1(_00600_),
    .A2(_01701_),
    .B1(_04105_),
    .B2(_04108_),
    .C(_04152_),
    .ZN(_04187_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _10079_ (.A1(_00847_),
    .A2(_01701_),
    .B(_01103_),
    .ZN(_04188_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10080_ (.A1(_04187_),
    .A2(_04188_),
    .ZN(_04189_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10081_ (.A1(_04186_),
    .A2(_04189_),
    .Z(_04190_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _10082_ (.A1(_00600_),
    .A2(_01712_),
    .B1(_04097_),
    .B2(_04100_),
    .C(_04147_),
    .ZN(_04191_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _10083_ (.A1(_00847_),
    .A2(_01712_),
    .B(_01038_),
    .ZN(_04192_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10084_ (.A1(_04191_),
    .A2(_04192_),
    .ZN(_04193_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10085_ (.A1(_04186_),
    .A2(_04193_),
    .Z(_04194_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10086_ (.I(_03840_),
    .Z(_04195_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10087_ (.A1(_03972_),
    .A2(_04190_),
    .B1(_04194_),
    .B2(_04195_),
    .ZN(_04196_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _10088_ (.A1(_03975_),
    .A2(_04177_),
    .B1(_04196_),
    .B2(_00766_),
    .C(_00764_),
    .ZN(_04197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10089_ (.A1(_04116_),
    .A2(_04169_),
    .ZN(_04198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10090_ (.A1(_04170_),
    .A2(_04198_),
    .ZN(_04199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10091_ (.A1(_04166_),
    .A2(_04199_),
    .ZN(_04200_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10092_ (.A1(_04166_),
    .A2(_04199_),
    .ZN(_04201_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10093_ (.A1(_00764_),
    .A2(_04201_),
    .ZN(_04202_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10094_ (.A1(_04200_),
    .A2(_04202_),
    .B(_04070_),
    .ZN(_04203_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10095_ (.A1(_04124_),
    .A2(_04184_),
    .B1(_04197_),
    .B2(_04203_),
    .ZN(_04204_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10096_ (.A1(_02185_),
    .A2(_03922_),
    .B1(_04204_),
    .B2(_03982_),
    .ZN(_04205_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10097_ (.I(_03806_),
    .Z(_04206_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10098_ (.A1(_04165_),
    .A2(_04206_),
    .B(_04122_),
    .ZN(_04207_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10099_ (.A1(_04036_),
    .A2(_04205_),
    .B(_04207_),
    .ZN(_00302_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10100_ (.I(_03747_),
    .Z(_04208_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10101_ (.A1(net92),
    .A2(_01621_),
    .ZN(_04209_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10102_ (.I(_04209_),
    .Z(_04210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10103_ (.A1(_02183_),
    .A2(_01624_),
    .ZN(_04211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10104_ (.A1(_04211_),
    .A2(_04200_),
    .ZN(_04212_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10105_ (.A1(_04210_),
    .A2(_04212_),
    .ZN(_04213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10106_ (.I(\as2650.addr_buff[1] ),
    .Z(_04214_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10107_ (.I(_04214_),
    .Z(_04215_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _10108_ (.A1(_04186_),
    .A2(_04191_),
    .A3(_04192_),
    .ZN(_04216_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10109_ (.A1(_04215_),
    .A2(_04216_),
    .Z(_04217_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _10110_ (.A1(_04185_),
    .A2(_04187_),
    .A3(_04188_),
    .ZN(_04218_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10111_ (.A1(_04214_),
    .A2(_04218_),
    .Z(_04219_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _10112_ (.A1(_04103_),
    .A2(_04217_),
    .B1(_04219_),
    .B2(_04112_),
    .ZN(_04220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10113_ (.I(net39),
    .Z(_04221_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10114_ (.A1(net38),
    .A2(_04176_),
    .ZN(_04222_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10115_ (.A1(_04221_),
    .A2(_04222_),
    .Z(_04223_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10116_ (.A1(_03797_),
    .A2(_04220_),
    .B1(_04223_),
    .B2(_03873_),
    .C(_04158_),
    .ZN(_04224_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10117_ (.A1(_03947_),
    .A2(_04213_),
    .B(_04224_),
    .ZN(_04225_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10118_ (.I(_04126_),
    .Z(_04226_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10119_ (.I(_03693_),
    .Z(_04227_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10120_ (.I(_04227_),
    .Z(_04228_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10121_ (.A1(_04215_),
    .A2(_03770_),
    .B1(_03772_),
    .B2(_04221_),
    .C(_01231_),
    .ZN(_04229_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10122_ (.A1(_04228_),
    .A2(_04223_),
    .B(_04229_),
    .ZN(_04230_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10123_ (.A1(_02196_),
    .A2(_04226_),
    .B(_04230_),
    .ZN(_04231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10124_ (.A1(_04166_),
    .A2(_04171_),
    .ZN(_04232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10125_ (.A1(_04211_),
    .A2(_04232_),
    .ZN(_04233_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10126_ (.A1(_04210_),
    .A2(_04233_),
    .Z(_04234_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10127_ (.A1(_03760_),
    .A2(_04234_),
    .ZN(_04235_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10128_ (.A1(_04221_),
    .A2(_03757_),
    .B(_04139_),
    .C(_04235_),
    .ZN(_04236_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10129_ (.A1(_00719_),
    .A2(_04231_),
    .B(_04236_),
    .ZN(_04237_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10130_ (.A1(_02197_),
    .A2(_04075_),
    .B1(_04237_),
    .B2(_04142_),
    .ZN(_04238_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10131_ (.A1(_03979_),
    .A2(_04225_),
    .B1(_04238_),
    .B2(_04124_),
    .ZN(_04239_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10132_ (.I(_03981_),
    .Z(_04240_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10133_ (.A1(_02197_),
    .A2(_03987_),
    .B1(_04239_),
    .B2(_04240_),
    .ZN(_04241_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10134_ (.A1(_04221_),
    .A2(_04206_),
    .B(_04122_),
    .ZN(_04242_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10135_ (.A1(_04208_),
    .A2(_04241_),
    .B(_04242_),
    .ZN(_00303_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10136_ (.I(_00541_),
    .Z(_04243_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10137_ (.I(_04243_),
    .Z(_04244_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10138_ (.I(_03812_),
    .Z(_04245_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10139_ (.A1(net39),
    .A2(net38),
    .A3(_04176_),
    .ZN(_04246_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10140_ (.A1(net96),
    .A2(_04246_),
    .Z(_04247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10141_ (.A1(_04076_),
    .A2(_04247_),
    .ZN(_04248_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _10142_ (.I(\as2650.addr_buff[2] ),
    .ZN(_04249_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10143_ (.I(_04249_),
    .Z(_04250_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _10144_ (.I(net96),
    .ZN(_04251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10145_ (.I(_02748_),
    .Z(_04252_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10146_ (.A1(_04250_),
    .A2(_03824_),
    .B1(_03826_),
    .B2(_04251_),
    .C(_04252_),
    .ZN(_04253_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10147_ (.A1(_02203_),
    .A2(_04245_),
    .B1(_04248_),
    .B2(_04253_),
    .ZN(_04254_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10148_ (.A1(net66),
    .A2(_01621_),
    .Z(_04255_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _10149_ (.I(_04255_),
    .ZN(_04256_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10150_ (.A1(net92),
    .A2(_02182_),
    .B(_01622_),
    .ZN(_04257_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10151_ (.A1(_04232_),
    .A2(_04210_),
    .B(_04257_),
    .ZN(_04258_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10152_ (.A1(_04256_),
    .A2(_04258_),
    .Z(_04259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10153_ (.A1(_04082_),
    .A2(_04259_),
    .ZN(_04260_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10154_ (.A1(net96),
    .A2(_03903_),
    .B(_03763_),
    .C(_04260_),
    .ZN(_04261_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10155_ (.A1(_04244_),
    .A2(_04254_),
    .B(_04261_),
    .ZN(_04262_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10156_ (.A1(_02204_),
    .A2(_03928_),
    .B1(_04262_),
    .B2(_03912_),
    .C(_03857_),
    .ZN(_04263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10157_ (.A1(_02195_),
    .A2(_02851_),
    .ZN(_04264_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10158_ (.A1(_04211_),
    .A2(_04264_),
    .ZN(_04265_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10159_ (.A1(_04200_),
    .A2(_04210_),
    .ZN(_04266_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10160_ (.A1(_04265_),
    .A2(_04266_),
    .ZN(_04267_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10161_ (.A1(_04256_),
    .A2(_04267_),
    .Z(_04268_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10162_ (.A1(\as2650.addr_buff[0] ),
    .A2(\as2650.addr_buff[1] ),
    .A3(\as2650.addr_buff[2] ),
    .ZN(_04269_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _10163_ (.A1(_04191_),
    .A2(_04192_),
    .A3(_04269_),
    .ZN(_04270_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10164_ (.I(_04214_),
    .Z(_04271_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10165_ (.I(\as2650.addr_buff[2] ),
    .Z(_04272_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10166_ (.A1(_04271_),
    .A2(_04216_),
    .B(_04272_),
    .ZN(_04273_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10167_ (.A1(_04270_),
    .A2(_04273_),
    .B(_00636_),
    .ZN(_04274_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _10168_ (.A1(_04187_),
    .A2(_04188_),
    .A3(_04269_),
    .ZN(_04275_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10169_ (.A1(_04271_),
    .A2(_04218_),
    .B(_04272_),
    .ZN(_04276_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10170_ (.A1(_04275_),
    .A2(_04276_),
    .B(_03972_),
    .ZN(_04277_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10171_ (.A1(_04274_),
    .A2(_04277_),
    .ZN(_04278_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10172_ (.A1(_03783_),
    .A2(_04247_),
    .B1(_04278_),
    .B2(_03797_),
    .C(_04158_),
    .ZN(_04279_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _10173_ (.A1(_00866_),
    .A2(_04268_),
    .B(_04279_),
    .C(_04070_),
    .ZN(_04280_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10174_ (.A1(_04263_),
    .A2(_04280_),
    .B(_03865_),
    .ZN(_04281_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10175_ (.A1(_02204_),
    .A2(_03751_),
    .B(_04281_),
    .ZN(_04282_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10176_ (.I(_00845_),
    .Z(_04283_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10177_ (.A1(net96),
    .A2(_04206_),
    .B(_04283_),
    .ZN(_04284_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10178_ (.A1(_04208_),
    .A2(_04282_),
    .B(_04284_),
    .ZN(_00304_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10179_ (.A1(net91),
    .A2(_04096_),
    .ZN(_04285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10180_ (.A1(_02202_),
    .A2(_04146_),
    .ZN(_04286_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10181_ (.A1(_04256_),
    .A2(_04267_),
    .B(_04286_),
    .ZN(_04287_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10182_ (.A1(_04285_),
    .A2(_04287_),
    .ZN(_04288_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10183_ (.I(\as2650.addr_buff[3] ),
    .Z(_04289_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10184_ (.A1(_04289_),
    .A2(_04270_),
    .Z(_04290_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10185_ (.I(\as2650.addr_buff[3] ),
    .Z(_04291_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10186_ (.A1(_04291_),
    .A2(_04275_),
    .Z(_04292_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _10187_ (.A1(_04063_),
    .A2(_04290_),
    .B1(_04292_),
    .B2(_04112_),
    .ZN(_04293_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10188_ (.A1(_04251_),
    .A2(_04246_),
    .ZN(_04294_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10189_ (.A1(net41),
    .A2(_04294_),
    .Z(_04295_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10190_ (.I(_04295_),
    .ZN(_04296_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10191_ (.A1(_03892_),
    .A2(_04293_),
    .B1(_04296_),
    .B2(_03873_),
    .C(_04158_),
    .ZN(_04297_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10192_ (.A1(_03780_),
    .A2(_04288_),
    .B(_04297_),
    .ZN(_04298_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10193_ (.I(net41),
    .Z(_04299_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10194_ (.A1(_04289_),
    .A2(_03770_),
    .B1(_03825_),
    .B2(_04299_),
    .C(_01231_),
    .ZN(_04300_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10195_ (.A1(_04228_),
    .A2(_04296_),
    .B(_04300_),
    .ZN(_04301_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10196_ (.A1(_02209_),
    .A2(_04226_),
    .B(_04301_),
    .ZN(_04302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10197_ (.A1(_04255_),
    .A2(_04258_),
    .ZN(_04303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10198_ (.A1(_04286_),
    .A2(_04303_),
    .ZN(_04304_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10199_ (.A1(_04285_),
    .A2(_04304_),
    .Z(_04305_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10200_ (.A1(_03760_),
    .A2(_04305_),
    .ZN(_04306_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10201_ (.A1(_04299_),
    .A2(_03757_),
    .B(_04139_),
    .C(_04306_),
    .ZN(_04307_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10202_ (.A1(_00719_),
    .A2(_04302_),
    .B(_04307_),
    .ZN(_04308_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10203_ (.A1(_02210_),
    .A2(_04075_),
    .B1(_04308_),
    .B2(_04142_),
    .ZN(_04309_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10204_ (.A1(_03979_),
    .A2(_04298_),
    .B1(_04309_),
    .B2(_04124_),
    .ZN(_04310_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10205_ (.A1(_02210_),
    .A2(_03987_),
    .B1(_04310_),
    .B2(_04240_),
    .ZN(_04311_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10206_ (.A1(_04299_),
    .A2(_04206_),
    .B(_04283_),
    .ZN(_04312_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10207_ (.A1(_04208_),
    .A2(_04311_),
    .B(_04312_),
    .ZN(_00305_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10208_ (.A1(_04256_),
    .A2(_04285_),
    .ZN(_04313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10209_ (.A1(net91),
    .A2(_04146_),
    .ZN(_04314_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10210_ (.A1(_04286_),
    .A2(_04257_),
    .A3(_04314_),
    .ZN(_04315_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10211_ (.A1(_04266_),
    .A2(_04313_),
    .B(_04315_),
    .ZN(_04316_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10212_ (.A1(net68),
    .A2(_01623_),
    .Z(_04317_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10213_ (.A1(_04316_),
    .A2(_04317_),
    .ZN(_04318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10214_ (.I(\as2650.addr_buff[4] ),
    .Z(_04319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10215_ (.A1(_04291_),
    .A2(_04275_),
    .ZN(_04320_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10216_ (.A1(_04319_),
    .A2(_04320_),
    .ZN(_04321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10217_ (.A1(_04291_),
    .A2(_04270_),
    .ZN(_04322_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10218_ (.A1(\as2650.addr_buff[4] ),
    .A2(_04322_),
    .ZN(_04323_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _10219_ (.A1(_04112_),
    .A2(_04321_),
    .B1(_04323_),
    .B2(_04063_),
    .ZN(_04324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10220_ (.A1(_04299_),
    .A2(_04294_),
    .ZN(_04325_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10221_ (.A1(net95),
    .A2(_04325_),
    .Z(_04326_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10222_ (.A1(_03892_),
    .A2(_04324_),
    .B1(_04326_),
    .B2(_03873_),
    .C(_00865_),
    .ZN(_04327_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10223_ (.A1(_03780_),
    .A2(_04318_),
    .B(_04327_),
    .ZN(_04328_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10224_ (.A1(net95),
    .A2(_04019_),
    .ZN(_04329_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10225_ (.A1(_04319_),
    .A2(_04020_),
    .B(_03825_),
    .ZN(_04330_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10226_ (.I(_02515_),
    .Z(_04331_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _10227_ (.A1(_00742_),
    .A2(_04326_),
    .B1(_04329_),
    .B2(_04330_),
    .C(_04331_),
    .ZN(_04332_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10228_ (.A1(_02216_),
    .A2(_04226_),
    .B(_04332_),
    .ZN(_04333_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10229_ (.A1(_04232_),
    .A2(_04209_),
    .ZN(_04334_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10230_ (.A1(_04334_),
    .A2(_04313_),
    .B(_04315_),
    .ZN(_04335_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10231_ (.A1(_04317_),
    .A2(_04335_),
    .ZN(_04336_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10232_ (.A1(_03903_),
    .A2(_04336_),
    .ZN(_04337_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10233_ (.A1(net95),
    .A2(_04038_),
    .B(_04139_),
    .ZN(_04338_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10234_ (.A1(_04125_),
    .A2(_04333_),
    .B1(_04337_),
    .B2(_04338_),
    .ZN(_04339_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10235_ (.A1(_02217_),
    .A2(_04075_),
    .B1(_04339_),
    .B2(_04142_),
    .ZN(_04340_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10236_ (.A1(_03979_),
    .A2(_04328_),
    .B1(_04340_),
    .B2(_00827_),
    .ZN(_04341_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10237_ (.A1(_02217_),
    .A2(_03987_),
    .B1(_04341_),
    .B2(_04240_),
    .ZN(_04342_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10238_ (.A1(net95),
    .A2(_03747_),
    .B(_04283_),
    .ZN(_04343_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10239_ (.A1(_04208_),
    .A2(_04342_),
    .B(_04343_),
    .ZN(_00306_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _10240_ (.A1(_02535_),
    .A2(_02540_),
    .B(_02541_),
    .C(_02493_),
    .ZN(_04344_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10241_ (.A1(_03707_),
    .A2(_03715_),
    .A3(_04344_),
    .ZN(_04345_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _10242_ (.A1(_02532_),
    .A2(_02533_),
    .A3(_03717_),
    .ZN(_04346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10243_ (.A1(_00608_),
    .A2(_00617_),
    .ZN(_04347_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10244_ (.A1(_03756_),
    .A2(_00609_),
    .B(_04347_),
    .ZN(_04348_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10245_ (.I(_03696_),
    .ZN(_04349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10246_ (.A1(_04349_),
    .A2(_03711_),
    .ZN(_04350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10247_ (.A1(_03732_),
    .A2(_03733_),
    .ZN(_04351_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10248_ (.A1(_03721_),
    .A2(_04348_),
    .B(_04350_),
    .C(_04351_),
    .ZN(_04352_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _10249_ (.A1(_00638_),
    .A2(_00651_),
    .A3(_00916_),
    .A4(_03728_),
    .ZN(_04353_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10250_ (.A1(_00770_),
    .A2(_04353_),
    .ZN(_04354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10251_ (.A1(_00473_),
    .A2(_00544_),
    .ZN(_04355_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10252_ (.A1(_03690_),
    .A2(_04355_),
    .B(_03742_),
    .C(_02501_),
    .ZN(_04356_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10253_ (.A1(_00626_),
    .A2(_00855_),
    .A3(_03720_),
    .ZN(_04357_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10254_ (.A1(_04019_),
    .A2(_00885_),
    .A3(_00658_),
    .A4(_04357_),
    .ZN(_04358_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10255_ (.A1(_03904_),
    .A2(_00717_),
    .ZN(_04359_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10256_ (.A1(_02335_),
    .A2(_02333_),
    .A3(_04359_),
    .ZN(_04360_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10257_ (.A1(_03613_),
    .A2(_03727_),
    .A3(_04358_),
    .A4(_04360_),
    .ZN(_04361_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10258_ (.A1(_04354_),
    .A2(_04356_),
    .A3(_04361_),
    .ZN(_04362_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10259_ (.A1(_04346_),
    .A2(_04352_),
    .A3(_04362_),
    .ZN(_04363_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _10260_ (.A1(_03706_),
    .A2(_04345_),
    .A3(_04363_),
    .Z(_04364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10261_ (.I(_03911_),
    .Z(_04365_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10262_ (.I(_00791_),
    .Z(_04366_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10263_ (.I(_04366_),
    .Z(_04367_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10264_ (.I(_04367_),
    .Z(_04368_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10265_ (.A1(net89),
    .A2(_04368_),
    .ZN(_04369_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10266_ (.A1(_03927_),
    .A2(_00503_),
    .ZN(_04370_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10267_ (.A1(_02903_),
    .A2(_04369_),
    .B(_04370_),
    .ZN(_04371_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10268_ (.I(_00739_),
    .Z(_04372_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10269_ (.A1(net28),
    .A2(_04372_),
    .A3(_04017_),
    .ZN(_04373_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10270_ (.A1(net28),
    .A2(_00592_),
    .B(_00654_),
    .C(_03800_),
    .ZN(_04374_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10271_ (.A1(_04365_),
    .A2(_04371_),
    .B(_04373_),
    .C(_04374_),
    .ZN(_04375_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10272_ (.A1(_03917_),
    .A2(_04375_),
    .B(_04364_),
    .ZN(_04376_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10273_ (.A1(net89),
    .A2(_04364_),
    .B(_04376_),
    .C(_03689_),
    .ZN(_00307_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10274_ (.A1(_00782_),
    .A2(_00893_),
    .A3(_00726_),
    .ZN(_04377_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10275_ (.A1(_00968_),
    .A2(_00690_),
    .ZN(_04378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10276_ (.A1(_04378_),
    .A2(_03733_),
    .ZN(_04379_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _10277_ (.A1(_00799_),
    .A2(_00738_),
    .A3(_00491_),
    .A4(_02334_),
    .Z(_04380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10278_ (.A1(_00738_),
    .A2(_00708_),
    .ZN(_04381_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _10279_ (.A1(_00518_),
    .A2(_04381_),
    .A3(_00702_),
    .A4(_03740_),
    .ZN(_04382_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10280_ (.A1(_04379_),
    .A2(_04380_),
    .A3(_04382_),
    .ZN(_04383_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _10281_ (.A1(_00679_),
    .A2(_00545_),
    .A3(_00732_),
    .A4(_04016_),
    .ZN(_04384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10282_ (.A1(_00738_),
    .A2(_00702_),
    .ZN(_04385_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10283_ (.A1(_00786_),
    .A2(_00695_),
    .A3(_03728_),
    .ZN(_04386_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _10284_ (.A1(_04384_),
    .A2(_04385_),
    .A3(_04386_),
    .Z(_04387_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10285_ (.A1(_03731_),
    .A2(_03738_),
    .A3(_04383_),
    .A4(_04387_),
    .ZN(_04388_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _10286_ (.A1(_04377_),
    .A2(net83),
    .A3(_03726_),
    .A4(_04388_),
    .Z(_04389_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _10287_ (.A1(_00518_),
    .A2(_00659_),
    .A3(_00663_),
    .A4(_03740_),
    .ZN(_04390_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10288_ (.I(_04390_),
    .ZN(_04391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10289_ (.A1(_02739_),
    .A2(_02932_),
    .ZN(_04392_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _10290_ (.A1(_00838_),
    .A2(_00829_),
    .A3(_02506_),
    .A4(_04392_),
    .ZN(_04393_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10291_ (.A1(_04366_),
    .A2(_00492_),
    .A3(_03766_),
    .ZN(_04394_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _10292_ (.A1(_00782_),
    .A2(_00466_),
    .ZN(_04395_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10293_ (.A1(_04393_),
    .A2(_04394_),
    .B(_04395_),
    .ZN(_04396_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10294_ (.A1(_04391_),
    .A2(_04396_),
    .ZN(_04397_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _10295_ (.A1(_03706_),
    .A2(_03719_),
    .A3(_04389_),
    .A4(_04397_),
    .ZN(_04398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10296_ (.A1(_00783_),
    .A2(_00767_),
    .ZN(_04399_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10297_ (.I(_00710_),
    .Z(_04400_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10298_ (.A1(_00739_),
    .A2(_04400_),
    .ZN(_04401_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _10299_ (.A1(_00739_),
    .A2(_00647_),
    .A3(_03897_),
    .B1(_00721_),
    .B2(_04401_),
    .ZN(_04402_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10300_ (.I(_04243_),
    .Z(_04403_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10301_ (.A1(net94),
    .A2(_04402_),
    .B(_04403_),
    .ZN(_04404_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _10302_ (.A1(_00861_),
    .A2(_04359_),
    .A3(_04404_),
    .Z(_04405_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10303_ (.I(_00805_),
    .Z(_04406_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10304_ (.A1(net94),
    .A2(_04406_),
    .A3(_03669_),
    .ZN(_04407_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10305_ (.A1(net94),
    .A2(_00892_),
    .A3(_00857_),
    .A4(_03810_),
    .ZN(_04408_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _10306_ (.A1(_03729_),
    .A2(_04405_),
    .A3(_04407_),
    .A4(_04408_),
    .ZN(_04409_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10307_ (.A1(_04399_),
    .A2(_04409_),
    .B(_02548_),
    .ZN(_04410_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10308_ (.A1(net94),
    .A2(_04398_),
    .B(_04283_),
    .ZN(_04411_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10309_ (.A1(_04398_),
    .A2(_04410_),
    .B(_04411_),
    .ZN(_00308_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _10310_ (.I(_03109_),
    .ZN(_04412_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10311_ (.A1(_00829_),
    .A2(_00709_),
    .ZN(_04413_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10312_ (.A1(_00724_),
    .A2(_00701_),
    .B1(_04413_),
    .B2(_03835_),
    .ZN(_04414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10313_ (.A1(_00609_),
    .A2(_03723_),
    .ZN(_04415_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10314_ (.A1(_00917_),
    .A2(_01056_),
    .ZN(_04416_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _10315_ (.I(_04416_),
    .ZN(_04417_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _10316_ (.A1(_00798_),
    .A2(_01802_),
    .ZN(_04418_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _10317_ (.A1(_00541_),
    .A2(_00800_),
    .A3(_04418_),
    .A4(_03655_),
    .ZN(_04419_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10318_ (.I(_01033_),
    .Z(_04420_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _10319_ (.A1(_00844_),
    .A2(_00654_),
    .B(_01018_),
    .C(_04420_),
    .ZN(_04421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10320_ (.A1(_02762_),
    .A2(_04421_),
    .ZN(_04422_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _10321_ (.A1(_03660_),
    .A2(_03676_),
    .A3(_04419_),
    .A4(_04422_),
    .ZN(_04423_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _10322_ (.A1(_03671_),
    .A2(_04415_),
    .B1(_04417_),
    .B2(_03914_),
    .C(_04423_),
    .ZN(_04424_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _10323_ (.I(_03898_),
    .Z(_04425_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10324_ (.A1(_00511_),
    .A2(_00786_),
    .A3(_00663_),
    .ZN(_04426_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10325_ (.A1(_04425_),
    .A2(_04385_),
    .A3(_04426_),
    .ZN(_04427_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _10326_ (.A1(_00627_),
    .A2(_00733_),
    .A3(_04016_),
    .A4(_04427_),
    .ZN(_04428_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10327_ (.A1(_00536_),
    .A2(_04414_),
    .B(_04424_),
    .C(_04428_),
    .ZN(_04429_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10328_ (.I(_04429_),
    .Z(_04430_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10329_ (.I(_04430_),
    .Z(_04431_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10330_ (.I(_04429_),
    .Z(_04432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10331_ (.A1(_04179_),
    .A2(_04432_),
    .ZN(_04433_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10332_ (.A1(_04412_),
    .A2(_04431_),
    .B(_04433_),
    .ZN(_00309_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10333_ (.I(_04429_),
    .Z(_04434_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10334_ (.A1(_04271_),
    .A2(_04434_),
    .ZN(_04435_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10335_ (.A1(_03886_),
    .A2(_04431_),
    .B(_04435_),
    .ZN(_00310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10336_ (.A1(_04272_),
    .A2(_04434_),
    .ZN(_04436_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10337_ (.A1(_03884_),
    .A2(_04431_),
    .B(_04436_),
    .ZN(_00311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10338_ (.A1(_04289_),
    .A2(_04434_),
    .ZN(_04437_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10339_ (.A1(_03951_),
    .A2(_04431_),
    .B(_04437_),
    .ZN(_00312_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10340_ (.I(_04319_),
    .Z(_04438_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10341_ (.A1(_04438_),
    .A2(_04434_),
    .ZN(_04439_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10342_ (.A1(_04003_),
    .A2(_04432_),
    .B(_04439_),
    .ZN(_00313_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _10343_ (.I(_01036_),
    .Z(_04440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10344_ (.A1(_04440_),
    .A2(_04430_),
    .ZN(_04441_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10345_ (.A1(_03203_),
    .A2(_04432_),
    .B(_04441_),
    .ZN(_00314_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10346_ (.I(_02854_),
    .Z(_04442_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 _10347_ (.I(_01035_),
    .Z(_04443_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10348_ (.I0(_04442_),
    .I1(_04443_),
    .S(_04430_),
    .Z(_04444_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10349_ (.I(_04444_),
    .Z(_00315_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10350_ (.A1(_00632_),
    .A2(_04430_),
    .ZN(_04445_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10351_ (.A1(_04038_),
    .A2(_04432_),
    .B(_04445_),
    .ZN(_00316_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10352_ (.A1(\as2650.last_intr ),
    .A2(_04033_),
    .ZN(_04446_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10353_ (.A1(_00689_),
    .A2(_02548_),
    .B(_04446_),
    .C(_03689_),
    .ZN(_00317_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10354_ (.I(_00914_),
    .Z(_04447_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10355_ (.A1(_04447_),
    .A2(_02332_),
    .B(_02537_),
    .C(_03689_),
    .ZN(_00318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10356_ (.A1(_03725_),
    .A2(_03742_),
    .ZN(_04448_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _10357_ (.A1(_00596_),
    .A2(_03721_),
    .B(_04448_),
    .ZN(_04449_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10358_ (.A1(_00624_),
    .A2(_03703_),
    .B1(_02536_),
    .B2(_02490_),
    .ZN(_04450_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10359_ (.A1(_04378_),
    .A2(_03732_),
    .A3(_04450_),
    .ZN(_04451_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10360_ (.A1(_03739_),
    .A2(_04451_),
    .ZN(_04452_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10361_ (.I(_03785_),
    .Z(_04453_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10362_ (.A1(_04453_),
    .A2(_00638_),
    .A3(_03721_),
    .ZN(_04454_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _10363_ (.A1(_00765_),
    .A2(_00756_),
    .A3(_00917_),
    .A4(_03729_),
    .ZN(_04455_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _10364_ (.A1(_04449_),
    .A2(_04452_),
    .A3(_04454_),
    .A4(_04455_),
    .ZN(_04456_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _10365_ (.A1(_04440_),
    .A2(_03917_),
    .B(_04456_),
    .ZN(_04457_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10366_ (.I(_03688_),
    .Z(_04458_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10367_ (.A1(_01193_),
    .A2(_04456_),
    .B(_04457_),
    .C(_04458_),
    .ZN(_00319_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _10368_ (.A1(_04443_),
    .A2(_03917_),
    .B(_04456_),
    .ZN(_04459_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10369_ (.A1(_01048_),
    .A2(_04456_),
    .B(_04459_),
    .C(_04458_),
    .ZN(_00320_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10370_ (.A1(_00792_),
    .A2(_02856_),
    .ZN(_04460_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10371_ (.A1(_01829_),
    .A2(_03762_),
    .B(_04460_),
    .ZN(_04461_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10372_ (.A1(_00902_),
    .A2(_00961_),
    .B(_00816_),
    .C(_01117_),
    .ZN(_04462_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10373_ (.A1(_02768_),
    .A2(_04462_),
    .B(_02335_),
    .ZN(_04463_));
 gf180mcu_fd_sc_mcu7t5v0__or3_2 _10374_ (.A1(_00894_),
    .A2(_01015_),
    .A3(_04463_),
    .Z(_04464_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10375_ (.I(_04464_),
    .Z(_04465_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10376_ (.I0(_04461_),
    .I1(_01099_),
    .S(_04465_),
    .Z(_04466_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10377_ (.I(_04466_),
    .Z(_00321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10378_ (.A1(_02560_),
    .A2(_03841_),
    .ZN(_04467_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10379_ (.I(_03832_),
    .Z(_04468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10380_ (.A1(_01850_),
    .A2(_04468_),
    .ZN(_04469_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _10381_ (.A1(_04467_),
    .A2(_04469_),
    .ZN(_04470_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10382_ (.I0(_04470_),
    .I1(\as2650.holding_reg[1] ),
    .S(_04465_),
    .Z(_04471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10383_ (.I(_04471_),
    .Z(_00322_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10384_ (.I(_04464_),
    .Z(_04472_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10385_ (.I(_00792_),
    .Z(_04473_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10386_ (.I(_04473_),
    .Z(_04474_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10387_ (.A1(_04474_),
    .A2(_03884_),
    .ZN(_04475_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _10388_ (.A1(_02067_),
    .A2(_00796_),
    .B(_04475_),
    .ZN(_04476_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10389_ (.I(_04464_),
    .Z(_04477_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10390_ (.A1(\as2650.holding_reg[2] ),
    .A2(_04477_),
    .ZN(_04478_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10391_ (.A1(_04472_),
    .A2(_04476_),
    .B(_04478_),
    .ZN(_00323_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10392_ (.A1(_00794_),
    .A2(_03951_),
    .ZN(_04479_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _10393_ (.A1(_02098_),
    .A2(_00796_),
    .B(_04479_),
    .ZN(_04480_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10394_ (.A1(\as2650.holding_reg[3] ),
    .A2(_04477_),
    .ZN(_04481_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10395_ (.A1(_04472_),
    .A2(_04480_),
    .B(_04481_),
    .ZN(_00324_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10396_ (.A1(_00537_),
    .A2(_04003_),
    .ZN(_04482_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10397_ (.A1(_03622_),
    .A2(_00796_),
    .B(_04482_),
    .ZN(_04483_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10398_ (.A1(\as2650.holding_reg[4] ),
    .A2(_04477_),
    .ZN(_04484_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10399_ (.A1(_04472_),
    .A2(_04483_),
    .B(_04484_),
    .ZN(_00325_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10400_ (.I(_04366_),
    .Z(_04485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10401_ (.A1(_01899_),
    .A2(_00583_),
    .ZN(_04486_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10402_ (.A1(_04485_),
    .A2(_04045_),
    .B(_04486_),
    .ZN(_04487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10403_ (.A1(\as2650.holding_reg[5] ),
    .A2(_04465_),
    .ZN(_04488_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10404_ (.A1(_04477_),
    .A2(_04487_),
    .B(_04488_),
    .ZN(_00326_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10405_ (.I(_03927_),
    .Z(_04489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10406_ (.A1(_02562_),
    .A2(_04442_),
    .ZN(_04490_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10407_ (.A1(_03625_),
    .A2(_04489_),
    .B(_04490_),
    .ZN(_04491_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10408_ (.I0(_04491_),
    .I1(\as2650.holding_reg[6] ),
    .S(_04464_),
    .Z(_04492_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10409_ (.I(_04492_),
    .Z(_00327_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10410_ (.I(\as2650.holding_reg[7] ),
    .ZN(_04493_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10411_ (.A1(_04489_),
    .A2(_00852_),
    .B(_04465_),
    .ZN(_04494_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10412_ (.A1(_04493_),
    .A2(_04472_),
    .B1(_04494_),
    .B2(_02345_),
    .ZN(_00328_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _10413_ (.I(_00838_),
    .Z(_04495_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _10414_ (.A1(_04495_),
    .A2(_00853_),
    .A3(_00857_),
    .A4(_04392_),
    .ZN(_04496_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10415_ (.A1(_00783_),
    .A2(_04496_),
    .B(_00668_),
    .ZN(_04497_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _10416_ (.I(_04497_),
    .Z(_04498_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10417_ (.I(_04497_),
    .Z(_04499_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _10418_ (.A1(_00784_),
    .A2(_02857_),
    .B(_04395_),
    .C(_04499_),
    .ZN(_04500_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10419_ (.A1(_05733_),
    .A2(_04498_),
    .B(_04500_),
    .ZN(_00329_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _10420_ (.I(_02858_),
    .Z(_04501_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _10421_ (.A1(_00784_),
    .A2(_04501_),
    .B(_04395_),
    .C(_04499_),
    .ZN(_04502_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10422_ (.A1(_05725_),
    .A2(_04498_),
    .B(_04502_),
    .ZN(_00330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _10423_ (.I(_02860_),
    .Z(_04503_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10424_ (.A1(_04503_),
    .A2(_00802_),
    .B1(_04498_),
    .B2(_00831_),
    .ZN(_04504_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10425_ (.I(_04504_),
    .ZN(_00331_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _10426_ (.A1(_02555_),
    .A2(_00854_),
    .B(_00668_),
    .C(_00783_),
    .ZN(_04505_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _10427_ (.A1(_00784_),
    .A2(_02555_),
    .B(_04395_),
    .C(_04499_),
    .ZN(_04506_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _10428_ (.A1(_01108_),
    .A2(_04505_),
    .B(_04506_),
    .ZN(_00332_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10429_ (.I(_00801_),
    .Z(_04507_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10430_ (.A1(_04442_),
    .A2(_04507_),
    .B1(_04498_),
    .B2(_01601_),
    .ZN(_04508_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10431_ (.I(_04508_),
    .ZN(_00333_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10432_ (.A1(_00852_),
    .A2(_04507_),
    .B1(_04499_),
    .B2(_01180_),
    .ZN(_04509_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10433_ (.I(_04509_),
    .ZN(_00334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10434_ (.A1(_00691_),
    .A2(_03736_),
    .ZN(_04510_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10435_ (.A1(_00624_),
    .A2(_00823_),
    .A3(_03703_),
    .ZN(_04511_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10436_ (.A1(_04510_),
    .A2(_04511_),
    .B(_00773_),
    .ZN(_00335_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10437_ (.A1(_00760_),
    .A2(_03735_),
    .ZN(_04512_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10438_ (.A1(_02520_),
    .A2(_04512_),
    .ZN(_04513_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _10439_ (.A1(_00781_),
    .A2(_00758_),
    .A3(_04384_),
    .A4(_04426_),
    .ZN(_04514_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _10440_ (.A1(_02538_),
    .A2(_03708_),
    .A3(_04514_),
    .ZN(_04515_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _10441_ (.A1(_04346_),
    .A2(_04449_),
    .A3(_04513_),
    .A4(_04515_),
    .ZN(_04516_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10442_ (.A1(_03710_),
    .A2(_04390_),
    .ZN(_04517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10443_ (.A1(_03613_),
    .A2(_03732_),
    .ZN(_04518_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _10444_ (.A1(_00517_),
    .A2(_00721_),
    .A3(_03896_),
    .A4(_04418_),
    .ZN(_04519_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10445_ (.A1(_02523_),
    .A2(_04510_),
    .ZN(_04520_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _10446_ (.A1(_04382_),
    .A2(_04518_),
    .A3(_04519_),
    .A4(_04520_),
    .ZN(_04521_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _10447_ (.A1(_04353_),
    .A2(_04387_),
    .A3(_04517_),
    .A4(_04521_),
    .ZN(_04522_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _10448_ (.A1(_02504_),
    .A2(_04345_),
    .A3(_04516_),
    .A4(_04522_),
    .ZN(_04523_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10449_ (.I(_04523_),
    .ZN(_04524_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10450_ (.I(_04524_),
    .Z(_04525_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10451_ (.I(_04525_),
    .Z(_04526_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10452_ (.A1(_03914_),
    .A2(_00968_),
    .ZN(_04527_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10453_ (.I(_04527_),
    .Z(_04528_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10454_ (.I(_03923_),
    .Z(_04529_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10455_ (.I(_00583_),
    .Z(_04530_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10456_ (.A1(_01836_),
    .A2(net84),
    .ZN(_04531_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10457_ (.A1(_00626_),
    .A2(_01601_),
    .ZN(_04532_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10458_ (.A1(_01835_),
    .A2(_00828_),
    .ZN(_04533_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10459_ (.A1(_03752_),
    .A2(_00480_),
    .ZN(_04534_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10460_ (.A1(_04533_),
    .A2(_04534_),
    .ZN(_04535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10461_ (.A1(net84),
    .A2(_04535_),
    .ZN(_04536_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10462_ (.A1(_04532_),
    .A2(_04536_),
    .ZN(_04537_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10463_ (.A1(_00458_),
    .A2(_04535_),
    .ZN(_04538_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10464_ (.A1(_03765_),
    .A2(_00458_),
    .B(_04538_),
    .ZN(_04539_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10465_ (.A1(_04531_),
    .A2(_04537_),
    .B1(_04539_),
    .B2(_04532_),
    .ZN(_04540_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10466_ (.I(_04413_),
    .Z(_04541_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10467_ (.A1(_03765_),
    .A2(_03904_),
    .ZN(_04542_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10468_ (.A1(_04024_),
    .A2(_03758_),
    .B(_04542_),
    .ZN(_04543_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10469_ (.A1(_04541_),
    .A2(_04543_),
    .ZN(_04544_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10470_ (.A1(_04412_),
    .A2(_03827_),
    .ZN(_04545_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10471_ (.A1(_04186_),
    .A2(_03899_),
    .B(_00746_),
    .ZN(_04546_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10472_ (.A1(_04545_),
    .A2(_04546_),
    .B(_00793_),
    .C(_03767_),
    .ZN(_04547_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10473_ (.A1(_04530_),
    .A2(_04540_),
    .B1(_04544_),
    .B2(_04547_),
    .C(_00740_),
    .ZN(_04548_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10474_ (.I(_01231_),
    .Z(_04549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10475_ (.A1(_05832_),
    .A2(_04227_),
    .ZN(_04550_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10476_ (.A1(_02856_),
    .A2(_04550_),
    .B(_02516_),
    .ZN(_04551_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _10477_ (.A1(_03768_),
    .A2(_04550_),
    .B(_04551_),
    .ZN(_04552_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10478_ (.I(_00512_),
    .Z(_04553_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10479_ (.A1(_01836_),
    .A2(_04549_),
    .B(_04552_),
    .C(_04553_),
    .ZN(_04554_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _10480_ (.A1(_04244_),
    .A2(_04548_),
    .A3(_04554_),
    .ZN(_04555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10481_ (.A1(_00542_),
    .A2(_03777_),
    .ZN(_04556_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10482_ (.A1(_03927_),
    .A2(_04543_),
    .B(_04556_),
    .ZN(_04557_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10483_ (.I(_00682_),
    .Z(_04558_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10484_ (.I(_04558_),
    .Z(_04559_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10485_ (.I(_01948_),
    .Z(_04560_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10486_ (.I(_01809_),
    .Z(_04561_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10487_ (.I(_04561_),
    .Z(_04562_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10488_ (.I(_01952_),
    .Z(_04563_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10489_ (.I(_04563_),
    .Z(_04564_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10490_ (.A1(\as2650.stack[8][0] ),
    .A2(_04562_),
    .B1(_04564_),
    .B2(\as2650.stack[9][0] ),
    .ZN(_04565_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10491_ (.I(_01958_),
    .Z(_04566_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10492_ (.I(_01962_),
    .Z(_04567_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10493_ (.I(_04567_),
    .Z(_04568_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10494_ (.A1(\as2650.stack[11][0] ),
    .A2(_04566_),
    .B1(_04568_),
    .B2(\as2650.stack[10][0] ),
    .ZN(_04569_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10495_ (.A1(_04560_),
    .A2(_04565_),
    .A3(_04569_),
    .ZN(_04570_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10496_ (.I(_01969_),
    .Z(_04571_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10497_ (.A1(\as2650.stack[15][0] ),
    .A2(_04566_),
    .B1(_04568_),
    .B2(\as2650.stack[14][0] ),
    .ZN(_04572_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10498_ (.I(_04561_),
    .Z(_04573_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10499_ (.I(_04563_),
    .Z(_04574_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10500_ (.A1(\as2650.stack[12][0] ),
    .A2(_04573_),
    .B1(_04574_),
    .B2(\as2650.stack[13][0] ),
    .ZN(_04575_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10501_ (.A1(_04571_),
    .A2(_04572_),
    .A3(_04575_),
    .ZN(_04576_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10502_ (.A1(_04570_),
    .A2(_04576_),
    .ZN(_04577_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10503_ (.A1(\as2650.stack[0][0] ),
    .A2(_02820_),
    .B1(_02821_),
    .B2(\as2650.stack[1][0] ),
    .ZN(_04578_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10504_ (.A1(\as2650.stack[3][0] ),
    .A2(_02828_),
    .B1(_02829_),
    .B2(\as2650.stack[2][0] ),
    .ZN(_04579_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10505_ (.A1(_02819_),
    .A2(_04578_),
    .A3(_04579_),
    .ZN(_04580_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10506_ (.A1(\as2650.stack[7][0] ),
    .A2(_02837_),
    .B1(_02829_),
    .B2(\as2650.stack[6][0] ),
    .ZN(_04581_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10507_ (.A1(\as2650.stack[4][0] ),
    .A2(_02835_),
    .B1(_01954_),
    .B2(\as2650.stack[5][0] ),
    .ZN(_04582_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10508_ (.A1(_02827_),
    .A2(_04581_),
    .A3(_04582_),
    .ZN(_04583_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10509_ (.A1(_04580_),
    .A2(_04583_),
    .B(_01943_),
    .ZN(_04584_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _10510_ (.A1(_02818_),
    .A2(_04577_),
    .B(_04584_),
    .ZN(_04585_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10511_ (.A1(_04559_),
    .A2(_04585_),
    .ZN(_04586_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10512_ (.I(_02747_),
    .Z(_04587_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10513_ (.I(_04587_),
    .Z(_04588_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10514_ (.A1(_03753_),
    .A2(_04588_),
    .B(_03923_),
    .ZN(_04589_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _10515_ (.A1(_04529_),
    .A2(_04555_),
    .A3(_04557_),
    .B1(_04586_),
    .B2(_04589_),
    .ZN(_04590_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10516_ (.A1(_01791_),
    .A2(_04527_),
    .ZN(_04591_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10517_ (.I(_04524_),
    .Z(_04592_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10518_ (.A1(_04528_),
    .A2(_04590_),
    .B1(_04591_),
    .B2(_03753_),
    .C(_04592_),
    .ZN(_04593_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10519_ (.A1(_03753_),
    .A2(_04526_),
    .B(_04593_),
    .C(_04458_),
    .ZN(_00336_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10520_ (.A1(_01854_),
    .A2(_03765_),
    .Z(_04594_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10521_ (.I(_04587_),
    .Z(_04595_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10522_ (.I(_01809_),
    .Z(_04596_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10523_ (.I(_01952_),
    .Z(_04597_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10524_ (.A1(\as2650.stack[8][1] ),
    .A2(_04596_),
    .B1(_04597_),
    .B2(\as2650.stack[9][1] ),
    .ZN(_04598_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10525_ (.A1(\as2650.stack[11][1] ),
    .A2(_01958_),
    .B1(_02030_),
    .B2(\as2650.stack[10][1] ),
    .ZN(_04599_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10526_ (.A1(_01948_),
    .A2(_04598_),
    .A3(_04599_),
    .ZN(_04600_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10527_ (.A1(\as2650.stack[15][1] ),
    .A2(_01958_),
    .B1(_04567_),
    .B2(\as2650.stack[14][1] ),
    .ZN(_04601_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10528_ (.A1(\as2650.stack[12][1] ),
    .A2(_04596_),
    .B1(_04597_),
    .B2(\as2650.stack[13][1] ),
    .ZN(_04602_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10529_ (.A1(_01969_),
    .A2(_04601_),
    .A3(_04602_),
    .ZN(_04603_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10530_ (.A1(_04600_),
    .A2(_04603_),
    .ZN(_04604_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10531_ (.A1(\as2650.stack[0][1] ),
    .A2(_04561_),
    .B1(_04563_),
    .B2(\as2650.stack[1][1] ),
    .ZN(_04605_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10532_ (.A1(\as2650.stack[3][1] ),
    .A2(_02823_),
    .B1(_04567_),
    .B2(\as2650.stack[2][1] ),
    .ZN(_04606_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10533_ (.A1(_01947_),
    .A2(_04605_),
    .A3(_04606_),
    .ZN(_04607_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10534_ (.A1(\as2650.stack[7][1] ),
    .A2(_02823_),
    .B1(_01963_),
    .B2(\as2650.stack[6][1] ),
    .ZN(_04608_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10535_ (.A1(\as2650.stack[4][1] ),
    .A2(_04561_),
    .B1(_04563_),
    .B2(\as2650.stack[5][1] ),
    .ZN(_04609_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10536_ (.A1(_01969_),
    .A2(_04608_),
    .A3(_04609_),
    .ZN(_04610_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10537_ (.A1(_04607_),
    .A2(_04610_),
    .B(_01942_),
    .ZN(_04611_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _10538_ (.A1(_02817_),
    .A2(_04604_),
    .B(_04611_),
    .ZN(_04612_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10539_ (.A1(_04595_),
    .A2(_04612_),
    .ZN(_04613_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10540_ (.I(_04558_),
    .Z(_04614_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10541_ (.A1(_04614_),
    .A2(_04594_),
    .B(_03754_),
    .ZN(_04615_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10542_ (.I(_00473_),
    .Z(_04616_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10543_ (.A1(_01854_),
    .A2(_03904_),
    .ZN(_04617_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10544_ (.A1(_04024_),
    .A2(_03821_),
    .B(_04617_),
    .ZN(_04618_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10545_ (.A1(_04215_),
    .A2(_04227_),
    .B(_00895_),
    .ZN(_04619_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10546_ (.A1(_03886_),
    .A2(_03773_),
    .B(_04619_),
    .ZN(_04620_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10547_ (.A1(_04413_),
    .A2(_04618_),
    .B1(_04594_),
    .B2(_03924_),
    .C(_04620_),
    .ZN(_04621_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10548_ (.I(_00460_),
    .Z(_04622_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10549_ (.I(_04622_),
    .Z(_04623_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10550_ (.A1(_03809_),
    .A2(_01835_),
    .Z(_04624_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10551_ (.A1(_01853_),
    .A2(_04534_),
    .Z(_04625_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10552_ (.I(_00460_),
    .Z(_04626_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10553_ (.A1(_01855_),
    .A2(_04534_),
    .B(_04626_),
    .ZN(_04627_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10554_ (.A1(_04623_),
    .A2(_04624_),
    .B1(_04625_),
    .B2(_04627_),
    .ZN(_04628_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10555_ (.A1(_02549_),
    .A2(_04628_),
    .ZN(_04629_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10556_ (.A1(_00584_),
    .A2(_04621_),
    .B(_04629_),
    .ZN(_04630_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _10557_ (.I(_02748_),
    .Z(_04631_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10558_ (.I(_04631_),
    .Z(_04632_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10559_ (.A1(_01079_),
    .A2(_05832_),
    .ZN(_04633_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10560_ (.A1(_03885_),
    .A2(_05826_),
    .Z(_04634_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10561_ (.A1(_04633_),
    .A2(_04634_),
    .B(_04020_),
    .ZN(_04635_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _10562_ (.A1(_04633_),
    .A2(_04634_),
    .B(_04635_),
    .ZN(_04636_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10563_ (.A1(_02858_),
    .A2(_04076_),
    .B(_04636_),
    .ZN(_04637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10564_ (.A1(_04252_),
    .A2(_04594_),
    .ZN(_04638_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10565_ (.A1(_04632_),
    .A2(_04637_),
    .B(_04638_),
    .ZN(_04639_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10566_ (.I(_00582_),
    .Z(_04640_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10567_ (.A1(_04640_),
    .A2(_04624_),
    .ZN(_04641_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10568_ (.A1(_04367_),
    .A2(_04618_),
    .B(_04641_),
    .C(_04243_),
    .ZN(_04642_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10569_ (.A1(_03911_),
    .A2(_04642_),
    .ZN(_04643_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10570_ (.A1(_04616_),
    .A2(_04630_),
    .B1(_04639_),
    .B2(_04372_),
    .C(_04643_),
    .ZN(_04644_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10571_ (.A1(_04613_),
    .A2(_04615_),
    .B(_04644_),
    .ZN(_04645_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10572_ (.A1(_04591_),
    .A2(_04594_),
    .B1(_04645_),
    .B2(_04528_),
    .C(_04592_),
    .ZN(_04646_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _10573_ (.A1(_03809_),
    .A2(_04526_),
    .B(_04646_),
    .C(_04458_),
    .ZN(_00337_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10574_ (.I(_04591_),
    .Z(_04647_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10575_ (.A1(_01854_),
    .A2(_01835_),
    .ZN(_04648_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _10576_ (.A1(_01867_),
    .A2(_04648_),
    .ZN(_04649_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10577_ (.A1(\as2650.stack[8][2] ),
    .A2(_02961_),
    .B1(_02962_),
    .B2(\as2650.stack[9][2] ),
    .ZN(_04650_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10578_ (.A1(\as2650.stack[11][2] ),
    .A2(_02951_),
    .B1(_02957_),
    .B2(\as2650.stack[10][2] ),
    .ZN(_04651_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10579_ (.A1(_02834_),
    .A2(_04650_),
    .A3(_04651_),
    .ZN(_04652_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10580_ (.A1(\as2650.stack[15][2] ),
    .A2(_01979_),
    .B1(_02957_),
    .B2(\as2650.stack[14][2] ),
    .ZN(_04653_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10581_ (.A1(\as2650.stack[12][2] ),
    .A2(_02961_),
    .B1(_02962_),
    .B2(\as2650.stack[13][2] ),
    .ZN(_04654_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10582_ (.A1(_02950_),
    .A2(_04653_),
    .A3(_04654_),
    .ZN(_04655_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10583_ (.A1(_04652_),
    .A2(_04655_),
    .ZN(_04656_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10584_ (.A1(\as2650.stack[0][2] ),
    .A2(_02961_),
    .B1(_02962_),
    .B2(\as2650.stack[1][2] ),
    .ZN(_04657_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10585_ (.A1(\as2650.stack[3][2] ),
    .A2(_01979_),
    .B1(_02030_),
    .B2(\as2650.stack[2][2] ),
    .ZN(_04658_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10586_ (.A1(_01948_),
    .A2(_04657_),
    .A3(_04658_),
    .ZN(_04659_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10587_ (.A1(\as2650.stack[7][2] ),
    .A2(_01979_),
    .B1(_02030_),
    .B2(\as2650.stack[6][2] ),
    .ZN(_04660_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10588_ (.A1(\as2650.stack[4][2] ),
    .A2(_04596_),
    .B1(_04597_),
    .B2(\as2650.stack[5][2] ),
    .ZN(_04661_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10589_ (.A1(_02950_),
    .A2(_04660_),
    .A3(_04661_),
    .ZN(_04662_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10590_ (.A1(_04659_),
    .A2(_04662_),
    .B(_02817_),
    .ZN(_04663_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _10591_ (.A1(_01943_),
    .A2(_04656_),
    .B(_04663_),
    .ZN(_04664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10592_ (.A1(_02567_),
    .A2(_04664_),
    .ZN(_04665_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10593_ (.I(_04558_),
    .Z(_04666_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10594_ (.I(_04666_),
    .Z(_04667_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10595_ (.A1(_04667_),
    .A2(_04649_),
    .B(_03912_),
    .ZN(_04668_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10596_ (.I(_04485_),
    .Z(_04669_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10597_ (.I(_02932_),
    .Z(_04670_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10598_ (.A1(_01867_),
    .A2(_04670_),
    .ZN(_04671_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10599_ (.A1(_02941_),
    .A2(_03907_),
    .B(_04671_),
    .ZN(_04672_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _10600_ (.A1(_04250_),
    .A2(_00927_),
    .B(_03900_),
    .C(_00747_),
    .ZN(_04673_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10601_ (.A1(_04541_),
    .A2(_04672_),
    .B1(_04649_),
    .B2(_04245_),
    .C(_04673_),
    .ZN(_04674_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10602_ (.A1(_01866_),
    .A2(_04648_),
    .Z(_04675_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10603_ (.A1(net57),
    .A2(_04625_),
    .Z(_04676_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10604_ (.A1(_01867_),
    .A2(_04625_),
    .B(_04626_),
    .ZN(_04677_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10605_ (.A1(_00461_),
    .A2(_04675_),
    .B1(_04676_),
    .B2(_04677_),
    .ZN(_04678_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10606_ (.A1(_04530_),
    .A2(_04678_),
    .ZN(_04679_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10607_ (.A1(_04669_),
    .A2(_04674_),
    .B(_04679_),
    .ZN(_04680_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10608_ (.I(_04331_),
    .Z(_04681_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10609_ (.I(_04331_),
    .Z(_04682_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10610_ (.A1(net10),
    .A2(_05819_),
    .Z(_04683_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10611_ (.A1(_01214_),
    .A2(_05826_),
    .ZN(_04684_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _10612_ (.A1(_04633_),
    .A2(_04634_),
    .B(_04684_),
    .ZN(_04685_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _10613_ (.A1(_04683_),
    .A2(_04685_),
    .Z(_04686_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _10614_ (.A1(_04683_),
    .A2(_04685_),
    .B(_03827_),
    .ZN(_04687_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10615_ (.A1(_02859_),
    .A2(_00927_),
    .ZN(_04688_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10616_ (.A1(_04686_),
    .A2(_04687_),
    .B(_04688_),
    .ZN(_04689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10617_ (.A1(_04682_),
    .A2(_04689_),
    .ZN(_04690_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10618_ (.A1(_04681_),
    .A2(_04675_),
    .B(_04690_),
    .ZN(_04691_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10619_ (.A1(_04485_),
    .A2(_04675_),
    .ZN(_04692_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10620_ (.A1(_03832_),
    .A2(_04672_),
    .B(_04692_),
    .C(_04243_),
    .ZN(_04693_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10621_ (.A1(_03754_),
    .A2(_04693_),
    .ZN(_04694_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10622_ (.A1(_04616_),
    .A2(_04680_),
    .B1(_04691_),
    .B2(_00741_),
    .C(_04694_),
    .ZN(_04695_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10623_ (.A1(_04665_),
    .A2(_04668_),
    .B(_04695_),
    .ZN(_04696_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10624_ (.I(_04528_),
    .Z(_04697_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10625_ (.I(_04524_),
    .Z(_04698_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10626_ (.I(_04698_),
    .Z(_04699_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10627_ (.A1(_04647_),
    .A2(_04649_),
    .B1(_04696_),
    .B2(_04697_),
    .C(_04699_),
    .ZN(_04700_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10628_ (.I(_04523_),
    .Z(_04701_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10629_ (.I(_00882_),
    .Z(_04702_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10630_ (.A1(_01868_),
    .A2(_04701_),
    .B(_04702_),
    .ZN(_04703_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10631_ (.A1(_04700_),
    .A2(_04703_),
    .ZN(_00338_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10632_ (.I(_04413_),
    .Z(_04704_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10633_ (.A1(_03921_),
    .A2(_00604_),
    .ZN(_04705_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10634_ (.A1(_02942_),
    .A2(_03937_),
    .B(_04705_),
    .ZN(_04706_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10635_ (.A1(_04704_),
    .A2(_04706_),
    .ZN(_04707_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _10636_ (.A1(_01866_),
    .A2(_01853_),
    .A3(_01834_),
    .ZN(_04708_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10637_ (.A1(_01877_),
    .A2(_04708_),
    .Z(_04709_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10638_ (.A1(_03951_),
    .A2(_00743_),
    .ZN(_04710_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _10639_ (.I(_04291_),
    .ZN(_04711_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10640_ (.A1(_04711_),
    .A2(_00928_),
    .B(_00748_),
    .ZN(_04712_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _10641_ (.A1(_03925_),
    .A2(_04709_),
    .B1(_04710_),
    .B2(_04712_),
    .C(_04368_),
    .ZN(_04713_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10642_ (.I(_00715_),
    .Z(_04714_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10643_ (.A1(_03921_),
    .A2(_04676_),
    .Z(_04715_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10644_ (.I(_04622_),
    .Z(_04716_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _10645_ (.I(_04709_),
    .ZN(_04717_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10646_ (.I(_04473_),
    .Z(_04718_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10647_ (.A1(_04716_),
    .A2(_04717_),
    .B(_04718_),
    .ZN(_04719_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10648_ (.A1(_00462_),
    .A2(_04715_),
    .B(_04719_),
    .ZN(_04720_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _10649_ (.A1(_04707_),
    .A2(_04713_),
    .B(_04714_),
    .C(_04720_),
    .ZN(_04721_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10650_ (.A1(_04669_),
    .A2(_04717_),
    .ZN(_04722_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10651_ (.A1(_04468_),
    .A2(_04706_),
    .B(_04722_),
    .C(_00543_),
    .ZN(_04723_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10652_ (.A1(_01327_),
    .A2(_05811_),
    .Z(_04724_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10653_ (.A1(_01264_),
    .A2(_05819_),
    .ZN(_04725_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10654_ (.I(_04725_),
    .ZN(_04726_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _10655_ (.A1(_04683_),
    .A2(_04685_),
    .B(_04726_),
    .ZN(_04727_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _10656_ (.A1(_04724_),
    .A2(_04727_),
    .ZN(_04728_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _10657_ (.A1(_04724_),
    .A2(_04727_),
    .ZN(_04729_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10658_ (.A1(_03897_),
    .A2(_04729_),
    .ZN(_04730_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10659_ (.A1(_02863_),
    .A2(_04425_),
    .ZN(_04731_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10660_ (.A1(_04728_),
    .A2(_04730_),
    .B(_04731_),
    .C(_04682_),
    .ZN(_04732_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10661_ (.A1(_04681_),
    .A2(_04709_),
    .B(_04732_),
    .C(_04372_),
    .ZN(_04733_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10662_ (.A1(_04365_),
    .A2(_04723_),
    .A3(_04733_),
    .ZN(_04734_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10663_ (.I(_04596_),
    .Z(_04735_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10664_ (.I(_04597_),
    .Z(_04736_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10665_ (.A1(\as2650.stack[8][3] ),
    .A2(_04735_),
    .B1(_04736_),
    .B2(\as2650.stack[9][3] ),
    .ZN(_04737_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10666_ (.A1(\as2650.stack[11][3] ),
    .A2(_01959_),
    .B1(_02031_),
    .B2(\as2650.stack[10][3] ),
    .ZN(_04738_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10667_ (.A1(_04560_),
    .A2(_04737_),
    .A3(_04738_),
    .ZN(_04739_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10668_ (.I(_04567_),
    .Z(_04740_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10669_ (.A1(\as2650.stack[15][3] ),
    .A2(_01959_),
    .B1(_04740_),
    .B2(\as2650.stack[14][3] ),
    .ZN(_04741_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10670_ (.A1(\as2650.stack[12][3] ),
    .A2(_04735_),
    .B1(_04736_),
    .B2(\as2650.stack[13][3] ),
    .ZN(_04742_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10671_ (.A1(_01970_),
    .A2(_04741_),
    .A3(_04742_),
    .ZN(_04743_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10672_ (.A1(_04739_),
    .A2(_04743_),
    .ZN(_04744_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10673_ (.A1(\as2650.stack[0][3] ),
    .A2(_04573_),
    .B1(_04574_),
    .B2(\as2650.stack[1][3] ),
    .ZN(_04745_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10674_ (.A1(\as2650.stack[3][3] ),
    .A2(_02824_),
    .B1(_04568_),
    .B2(\as2650.stack[2][3] ),
    .ZN(_04746_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10675_ (.A1(_02819_),
    .A2(_04745_),
    .A3(_04746_),
    .ZN(_04747_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10676_ (.A1(\as2650.stack[7][3] ),
    .A2(_02824_),
    .B1(_01964_),
    .B2(\as2650.stack[6][3] ),
    .ZN(_04748_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10677_ (.A1(\as2650.stack[4][3] ),
    .A2(_04573_),
    .B1(_04574_),
    .B2(\as2650.stack[5][3] ),
    .ZN(_04749_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10678_ (.A1(_04571_),
    .A2(_04748_),
    .A3(_04749_),
    .ZN(_04750_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10679_ (.A1(_04747_),
    .A2(_04750_),
    .B(_02946_),
    .ZN(_04751_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _10680_ (.A1(_02818_),
    .A2(_04744_),
    .B(_04751_),
    .ZN(_04752_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10681_ (.A1(_04588_),
    .A2(_04752_),
    .ZN(_04753_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10682_ (.A1(_02567_),
    .A2(_04717_),
    .B(_04753_),
    .C(_00877_),
    .ZN(_04754_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10683_ (.A1(_04721_),
    .A2(_04734_),
    .B(_04754_),
    .C(_04697_),
    .ZN(_04755_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10684_ (.A1(_04647_),
    .A2(_04709_),
    .B(_04699_),
    .ZN(_04756_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10685_ (.I(_00507_),
    .Z(_04757_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10686_ (.A1(_01877_),
    .A2(_04526_),
    .B1(_04755_),
    .B2(_04756_),
    .C(_04757_),
    .ZN(_00339_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10687_ (.I(_04525_),
    .Z(_04758_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10688_ (.A1(_03920_),
    .A2(_04676_),
    .Z(_04759_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10689_ (.A1(_04014_),
    .A2(_04759_),
    .ZN(_04760_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10690_ (.A1(_04015_),
    .A2(_04759_),
    .Z(_04761_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10691_ (.A1(_00462_),
    .A2(_04760_),
    .A3(_04761_),
    .ZN(_04762_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10692_ (.A1(_01877_),
    .A2(_04708_),
    .ZN(_04763_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10693_ (.A1(_04014_),
    .A2(_04763_),
    .Z(_04764_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10694_ (.A1(_00888_),
    .A2(_04764_),
    .B(_03663_),
    .ZN(_04765_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10695_ (.A1(_04015_),
    .A2(_03905_),
    .ZN(_04766_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10696_ (.A1(_00604_),
    .A2(_04026_),
    .B(_04766_),
    .ZN(_04767_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10697_ (.A1(_04319_),
    .A2(_04228_),
    .ZN(_04768_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10698_ (.A1(_02849_),
    .A2(_04049_),
    .B(_04400_),
    .ZN(_04769_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10699_ (.A1(_04768_),
    .A2(_04769_),
    .B(_02561_),
    .ZN(_04770_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10700_ (.A1(_03925_),
    .A2(_04764_),
    .B1(_04767_),
    .B2(_04704_),
    .C(_04770_),
    .ZN(_04771_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _10701_ (.A1(_04762_),
    .A2(_04765_),
    .B(_04771_),
    .C(_04714_),
    .ZN(_04772_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10702_ (.I(_04631_),
    .Z(_04773_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10703_ (.A1(_02849_),
    .A2(_04048_),
    .ZN(_04774_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10704_ (.A1(_01423_),
    .A2(_05801_),
    .Z(_04775_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10705_ (.A1(_02862_),
    .A2(_05811_),
    .ZN(_04776_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10706_ (.A1(_04724_),
    .A2(_04727_),
    .B(_04776_),
    .ZN(_04777_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10707_ (.A1(_04775_),
    .A2(_04777_),
    .ZN(_04778_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10708_ (.A1(_04775_),
    .A2(_04777_),
    .Z(_04779_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _10709_ (.A1(_03897_),
    .A2(_04778_),
    .A3(_04779_),
    .ZN(_04780_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10710_ (.A1(_04774_),
    .A2(_04780_),
    .B(_04773_),
    .ZN(_04781_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10711_ (.A1(_04773_),
    .A2(_04764_),
    .B(_04781_),
    .ZN(_04782_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10712_ (.A1(_01889_),
    .A2(_04763_),
    .Z(_04783_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10713_ (.A1(_04474_),
    .A2(_04783_),
    .ZN(_04784_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10714_ (.A1(_00537_),
    .A2(_04767_),
    .B(_04784_),
    .C(_04244_),
    .ZN(_04785_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10715_ (.A1(_00514_),
    .A2(_04782_),
    .B(_04785_),
    .C(_04365_),
    .ZN(_04786_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10716_ (.A1(\as2650.stack[8][4] ),
    .A2(_04562_),
    .B1(_04564_),
    .B2(\as2650.stack[9][4] ),
    .ZN(_04787_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10717_ (.A1(\as2650.stack[11][4] ),
    .A2(_01959_),
    .B1(_04740_),
    .B2(\as2650.stack[10][4] ),
    .ZN(_04788_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10718_ (.A1(_04560_),
    .A2(_04787_),
    .A3(_04788_),
    .ZN(_04789_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10719_ (.A1(\as2650.stack[15][4] ),
    .A2(_04566_),
    .B1(_04740_),
    .B2(\as2650.stack[14][4] ),
    .ZN(_04790_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10720_ (.A1(\as2650.stack[12][4] ),
    .A2(_04562_),
    .B1(_04564_),
    .B2(\as2650.stack[13][4] ),
    .ZN(_04791_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10721_ (.A1(_04571_),
    .A2(_04790_),
    .A3(_04791_),
    .ZN(_04792_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10722_ (.A1(_04789_),
    .A2(_04792_),
    .ZN(_04793_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10723_ (.A1(\as2650.stack[0][4] ),
    .A2(_02820_),
    .B1(_02821_),
    .B2(\as2650.stack[1][4] ),
    .ZN(_04794_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10724_ (.A1(\as2650.stack[3][4] ),
    .A2(_02828_),
    .B1(_01964_),
    .B2(\as2650.stack[2][4] ),
    .ZN(_04795_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10725_ (.A1(_02819_),
    .A2(_04794_),
    .A3(_04795_),
    .ZN(_04796_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10726_ (.A1(\as2650.stack[7][4] ),
    .A2(_02828_),
    .B1(_02829_),
    .B2(\as2650.stack[6][4] ),
    .ZN(_04797_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10727_ (.A1(\as2650.stack[4][4] ),
    .A2(_02835_),
    .B1(_01954_),
    .B2(\as2650.stack[5][4] ),
    .ZN(_04798_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10728_ (.A1(_02827_),
    .A2(_04797_),
    .A3(_04798_),
    .ZN(_04799_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10729_ (.A1(_04796_),
    .A2(_04799_),
    .B(_02946_),
    .ZN(_04800_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _10730_ (.A1(_02818_),
    .A2(_04793_),
    .B(_04800_),
    .ZN(_04801_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10731_ (.A1(_04588_),
    .A2(_04801_),
    .ZN(_04802_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10732_ (.A1(_02567_),
    .A2(_04783_),
    .B(_04802_),
    .C(_00877_),
    .ZN(_04803_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10733_ (.A1(_04772_),
    .A2(_04786_),
    .B(_04803_),
    .C(_04697_),
    .ZN(_04804_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10734_ (.A1(_04647_),
    .A2(_04764_),
    .B(_04699_),
    .ZN(_04805_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _10735_ (.I(_03688_),
    .Z(_04806_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10736_ (.A1(_01889_),
    .A2(_04758_),
    .B1(_04804_),
    .B2(_04805_),
    .C(_04806_),
    .ZN(_00340_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _10737_ (.A1(_01888_),
    .A2(_01876_),
    .A3(_04708_),
    .ZN(_04807_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10738_ (.A1(_01902_),
    .A2(_04807_),
    .Z(_04808_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10739_ (.I(_04808_),
    .Z(_04809_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10740_ (.A1(\as2650.stack[8][5] ),
    .A2(_04735_),
    .B1(_04736_),
    .B2(\as2650.stack[9][5] ),
    .ZN(_04810_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10741_ (.A1(\as2650.stack[11][5] ),
    .A2(_01980_),
    .B1(_02031_),
    .B2(\as2650.stack[10][5] ),
    .ZN(_04811_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10742_ (.A1(_01949_),
    .A2(_04810_),
    .A3(_04811_),
    .ZN(_04812_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10743_ (.A1(\as2650.stack[15][5] ),
    .A2(_01980_),
    .B1(_02031_),
    .B2(\as2650.stack[14][5] ),
    .ZN(_04813_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10744_ (.A1(\as2650.stack[12][5] ),
    .A2(_04735_),
    .B1(_04736_),
    .B2(\as2650.stack[13][5] ),
    .ZN(_04814_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10745_ (.A1(_01970_),
    .A2(_04813_),
    .A3(_04814_),
    .ZN(_04815_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10746_ (.A1(_04812_),
    .A2(_04815_),
    .ZN(_04816_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10747_ (.A1(\as2650.stack[0][5] ),
    .A2(_04562_),
    .B1(_04564_),
    .B2(\as2650.stack[1][5] ),
    .ZN(_04817_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10748_ (.A1(\as2650.stack[3][5] ),
    .A2(_04566_),
    .B1(_04740_),
    .B2(\as2650.stack[2][5] ),
    .ZN(_04818_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10749_ (.A1(_04560_),
    .A2(_04817_),
    .A3(_04818_),
    .ZN(_04819_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10750_ (.A1(\as2650.stack[7][5] ),
    .A2(_02824_),
    .B1(_04568_),
    .B2(\as2650.stack[6][5] ),
    .ZN(_04820_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10751_ (.A1(\as2650.stack[4][5] ),
    .A2(_04573_),
    .B1(_04574_),
    .B2(\as2650.stack[5][5] ),
    .ZN(_04821_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10752_ (.A1(_04571_),
    .A2(_04820_),
    .A3(_04821_),
    .ZN(_04822_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10753_ (.A1(_04819_),
    .A2(_04822_),
    .B(_02946_),
    .ZN(_04823_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _10754_ (.A1(_01944_),
    .A2(_04816_),
    .B(_04823_),
    .ZN(_04824_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10755_ (.A1(_04614_),
    .A2(_04824_),
    .ZN(_04825_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10756_ (.I(_00876_),
    .Z(_04826_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10757_ (.A1(_04588_),
    .A2(_04809_),
    .B(_04826_),
    .ZN(_04827_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10758_ (.I(_00513_),
    .Z(_04828_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10759_ (.A1(_02553_),
    .A2(_04425_),
    .ZN(_04829_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10760_ (.A1(_01535_),
    .A2(_05789_),
    .Z(_04830_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10761_ (.A1(_01424_),
    .A2(_05801_),
    .ZN(_04831_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _10762_ (.I(_04831_),
    .ZN(_04832_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10763_ (.A1(_04775_),
    .A2(_04777_),
    .B(_04832_),
    .ZN(_04833_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10764_ (.A1(_04830_),
    .A2(_04833_),
    .B(_00787_),
    .ZN(_04834_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10765_ (.A1(_04830_),
    .A2(_04833_),
    .B(_04834_),
    .ZN(_04835_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _10766_ (.A1(_04829_),
    .A2(_04835_),
    .B(_04631_),
    .ZN(_04836_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10767_ (.A1(_04549_),
    .A2(_04808_),
    .B(_04836_),
    .ZN(_04837_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10768_ (.A1(_01902_),
    .A2(_04760_),
    .Z(_04838_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10769_ (.A1(_00887_),
    .A2(_04808_),
    .ZN(_04839_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10770_ (.A1(_00887_),
    .A2(_04838_),
    .B(_04839_),
    .ZN(_04840_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10771_ (.A1(_00602_),
    .A2(_04042_),
    .ZN(_04841_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10772_ (.A1(_01903_),
    .A2(_00849_),
    .B(_04841_),
    .ZN(_04842_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10773_ (.A1(_01036_),
    .A2(_00661_),
    .ZN(_04843_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10774_ (.A1(_03203_),
    .A2(_03898_),
    .B(_04843_),
    .ZN(_04844_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10775_ (.A1(_03812_),
    .A2(_04808_),
    .B1(_04844_),
    .B2(_00895_),
    .C(_00792_),
    .ZN(_04845_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10776_ (.A1(_00859_),
    .A2(_04842_),
    .B(_04845_),
    .ZN(_04846_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10777_ (.A1(_03662_),
    .A2(_04840_),
    .B(_04846_),
    .C(_00513_),
    .ZN(_04847_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10778_ (.A1(_04828_),
    .A2(_04837_),
    .B(_04847_),
    .C(_00853_),
    .ZN(_04848_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10779_ (.A1(_00536_),
    .A2(_04809_),
    .ZN(_04849_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10780_ (.A1(_04718_),
    .A2(_04842_),
    .B(_04849_),
    .C(_00542_),
    .ZN(_04850_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10781_ (.A1(_03754_),
    .A2(_04848_),
    .A3(_04850_),
    .ZN(_04851_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10782_ (.A1(_04825_),
    .A2(_04827_),
    .B(_03679_),
    .C(_04851_),
    .ZN(_04852_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10783_ (.A1(_03680_),
    .A2(_04809_),
    .B(_04852_),
    .C(_00777_),
    .ZN(_04853_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10784_ (.I(_01791_),
    .Z(_04854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10785_ (.I(_04854_),
    .Z(_04855_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10786_ (.I(_02521_),
    .Z(_04856_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10787_ (.I(_04856_),
    .Z(_04857_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10788_ (.A1(\as2650.ivec[0] ),
    .A2(_04855_),
    .B1(_04857_),
    .B2(_04809_),
    .C(_04525_),
    .ZN(_04858_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10789_ (.A1(_04087_),
    .A2(_04758_),
    .B1(_04853_),
    .B2(_04858_),
    .C(_04806_),
    .ZN(_00341_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _10790_ (.I(_01912_),
    .ZN(_04859_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10791_ (.I(_04859_),
    .Z(_04860_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10792_ (.A1(_01902_),
    .A2(_04807_),
    .ZN(_04861_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10793_ (.A1(_04859_),
    .A2(_04861_),
    .Z(_04862_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10794_ (.I(_02516_),
    .Z(_04863_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10795_ (.A1(_01622_),
    .A2(_05857_),
    .Z(_04864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10796_ (.A1(_02552_),
    .A2(_05789_),
    .ZN(_04865_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10797_ (.A1(_04830_),
    .A2(_04833_),
    .B(_04865_),
    .ZN(_04866_));
 gf180mcu_fd_sc_mcu7t5v0__and2_2 _10798_ (.A1(_04864_),
    .A2(_04866_),
    .Z(_04867_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10799_ (.A1(_04864_),
    .A2(_04866_),
    .B(_03827_),
    .ZN(_04868_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10800_ (.A1(_02852_),
    .A2(_04425_),
    .ZN(_04869_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _10801_ (.A1(_04867_),
    .A2(_04868_),
    .B(_04869_),
    .ZN(_04870_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10802_ (.A1(_01912_),
    .A2(_01901_),
    .A3(_04807_),
    .ZN(_04871_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10803_ (.A1(_04860_),
    .A2(_04861_),
    .ZN(_04872_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10804_ (.A1(_04871_),
    .A2(_04872_),
    .ZN(_04873_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10805_ (.A1(_04331_),
    .A2(_04873_),
    .ZN(_04874_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10806_ (.A1(_04863_),
    .A2(_04870_),
    .B(_04874_),
    .ZN(_04875_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _10807_ (.A1(_01901_),
    .A2(_03988_),
    .A3(_04759_),
    .ZN(_04876_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10808_ (.A1(_04860_),
    .A2(_04876_),
    .Z(_04877_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10809_ (.A1(_04626_),
    .A2(_04877_),
    .ZN(_04878_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10810_ (.A1(_04623_),
    .A2(_04873_),
    .B(_04878_),
    .C(_04473_),
    .ZN(_04879_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10811_ (.A1(_00849_),
    .A2(_04091_),
    .ZN(_04880_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10812_ (.A1(_01913_),
    .A2(_04670_),
    .B(_04880_),
    .ZN(_04881_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10813_ (.A1(_04443_),
    .A2(_03898_),
    .ZN(_04882_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10814_ (.A1(_02851_),
    .A2(_00699_),
    .ZN(_04883_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10815_ (.A1(_04882_),
    .A2(_04883_),
    .ZN(_04884_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10816_ (.I(_00791_),
    .Z(_04885_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10817_ (.A1(_03812_),
    .A2(_04862_),
    .B1(_04884_),
    .B2(_00710_),
    .C(_04885_),
    .ZN(_04886_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10818_ (.A1(_00860_),
    .A2(_04881_),
    .B(_04886_),
    .ZN(_04887_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10819_ (.A1(_04553_),
    .A2(_04879_),
    .A3(_04887_),
    .ZN(_04888_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10820_ (.A1(_04828_),
    .A2(_04875_),
    .B(_04888_),
    .C(_00853_),
    .ZN(_04889_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10821_ (.I(_03762_),
    .Z(_04890_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10822_ (.A1(_04890_),
    .A2(_04862_),
    .ZN(_04891_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10823_ (.A1(_04669_),
    .A2(_04881_),
    .B(_04891_),
    .C(_04403_),
    .ZN(_04892_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10824_ (.A1(_00834_),
    .A2(_04889_),
    .A3(_04892_),
    .ZN(_04893_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10825_ (.A1(_04666_),
    .A2(_04873_),
    .ZN(_04894_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10826_ (.A1(_04614_),
    .A2(_02846_),
    .B(_04894_),
    .C(_04826_),
    .ZN(_04895_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10827_ (.A1(_00827_),
    .A2(_04893_),
    .A3(_04895_),
    .ZN(_04896_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10828_ (.A1(_03680_),
    .A2(_04862_),
    .B(_04896_),
    .C(_00777_),
    .ZN(_04897_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10829_ (.A1(\as2650.ivec[1] ),
    .A2(_04855_),
    .B1(_04857_),
    .B2(_04862_),
    .C(_04525_),
    .ZN(_04898_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10830_ (.A1(_04860_),
    .A2(_04758_),
    .B1(_04897_),
    .B2(_04898_),
    .C(_04806_),
    .ZN(_00342_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10831_ (.I(_04133_),
    .Z(_04899_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10832_ (.A1(_04899_),
    .A2(_04871_),
    .Z(_04900_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10833_ (.I(_04900_),
    .Z(_04901_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10834_ (.A1(_04899_),
    .A2(_03756_),
    .ZN(_04902_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10835_ (.A1(_03757_),
    .A2(_04137_),
    .B(_04902_),
    .ZN(_04903_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10836_ (.A1(_04019_),
    .A2(_04020_),
    .ZN(_04904_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10837_ (.A1(_03756_),
    .A2(_03773_),
    .B(_04904_),
    .ZN(_04905_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10838_ (.A1(_03924_),
    .A2(_04900_),
    .B1(_04905_),
    .B2(_04400_),
    .C(_00793_),
    .ZN(_04906_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10839_ (.A1(_00860_),
    .A2(_04903_),
    .B(_04906_),
    .ZN(_04907_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _10840_ (.A1(_04133_),
    .A2(_04859_),
    .A3(_04876_),
    .ZN(_04908_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10841_ (.A1(_04860_),
    .A2(_04876_),
    .ZN(_04909_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10842_ (.A1(net63),
    .A2(_04909_),
    .B(_00461_),
    .ZN(_04910_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10843_ (.A1(_00888_),
    .A2(_04900_),
    .ZN(_04911_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10844_ (.A1(_04908_),
    .A2(_04910_),
    .B(_04911_),
    .C(_04890_),
    .ZN(_04912_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10845_ (.A1(_04907_),
    .A2(_04912_),
    .B(_00715_),
    .ZN(_04913_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10846_ (.A1(_04530_),
    .A2(_04903_),
    .ZN(_04914_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _10847_ (.A1(_04368_),
    .A2(_04900_),
    .B(_04914_),
    .C(_04125_),
    .ZN(_04915_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10848_ (.A1(_03818_),
    .A2(_04049_),
    .ZN(_04916_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _10849_ (.A1(_01624_),
    .A2(_05857_),
    .B(_04867_),
    .ZN(_04917_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_2 _10850_ (.A1(_01705_),
    .A2(_05778_),
    .A3(_04917_),
    .Z(_04918_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10851_ (.A1(_04228_),
    .A2(_04918_),
    .ZN(_04919_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _10852_ (.A1(_04916_),
    .A2(_04919_),
    .B(_04549_),
    .ZN(_04920_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _10853_ (.A1(_04773_),
    .A2(_04901_),
    .B(_04920_),
    .C(_04828_),
    .ZN(_04921_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _10854_ (.A1(_04529_),
    .A2(_04913_),
    .A3(_04915_),
    .A4(_04921_),
    .ZN(_04922_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10855_ (.A1(_04595_),
    .A2(_04901_),
    .ZN(_04923_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10856_ (.A1(_04614_),
    .A2(_02966_),
    .B(_04826_),
    .ZN(_04924_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10857_ (.A1(_04923_),
    .A2(_04924_),
    .B(_00827_),
    .ZN(_04925_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _10858_ (.A1(_03680_),
    .A2(_04901_),
    .B1(_04922_),
    .B2(_04925_),
    .C(_03865_),
    .ZN(_04926_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10859_ (.A1(\as2650.ivec[2] ),
    .A2(_04855_),
    .B1(_04857_),
    .B2(_04901_),
    .C(_04592_),
    .ZN(_04927_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10860_ (.A1(_04899_),
    .A2(_04758_),
    .B1(_04926_),
    .B2(_04927_),
    .C(_04806_),
    .ZN(_00343_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _10861_ (.I(_04523_),
    .Z(_04928_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10862_ (.I(_03836_),
    .Z(_04929_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10863_ (.A1(_04899_),
    .A2(_04871_),
    .ZN(_04930_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_2 _10864_ (.A1(_02183_),
    .A2(_04930_),
    .ZN(_04931_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10865_ (.I(_04931_),
    .Z(_04932_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10866_ (.A1(_02184_),
    .A2(_04908_),
    .Z(_04933_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10867_ (.A1(_04716_),
    .A2(_04933_),
    .ZN(_04934_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10868_ (.A1(_04716_),
    .A2(_04932_),
    .B(_04934_),
    .C(_04890_),
    .ZN(_04935_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10869_ (.A1(_04670_),
    .A2(_04172_),
    .ZN(_04936_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10870_ (.A1(_02184_),
    .A2(_04670_),
    .Z(_04937_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10871_ (.A1(_04936_),
    .A2(_04937_),
    .ZN(_04938_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _10872_ (.A1(_04412_),
    .A2(_03899_),
    .B(_04180_),
    .C(_00746_),
    .ZN(_04939_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10873_ (.A1(_04485_),
    .A2(_04939_),
    .ZN(_04940_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _10874_ (.A1(_04226_),
    .A2(_04931_),
    .B1(_04938_),
    .B2(_00860_),
    .C(_04940_),
    .ZN(_04941_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10875_ (.A1(_04616_),
    .A2(_04935_),
    .A3(_04941_),
    .ZN(_04942_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10876_ (.A1(_02910_),
    .A2(_05778_),
    .ZN(_04943_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10877_ (.A1(_00601_),
    .A2(_05778_),
    .ZN(_04944_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _10878_ (.A1(_04943_),
    .A2(_04917_),
    .B(_04944_),
    .ZN(_04945_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10879_ (.A1(_04227_),
    .A2(_04945_),
    .Z(_04946_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10880_ (.A1(_04179_),
    .A2(_04946_),
    .Z(_04947_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10881_ (.A1(_04632_),
    .A2(_04932_),
    .ZN(_04948_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10882_ (.A1(_04773_),
    .A2(_04947_),
    .B(_04948_),
    .C(_04372_),
    .ZN(_04949_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10883_ (.A1(_04890_),
    .A2(_04931_),
    .B(_00718_),
    .ZN(_04950_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _10884_ (.A1(_00794_),
    .A2(_04936_),
    .A3(_04937_),
    .B(_04950_),
    .ZN(_04951_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _10885_ (.A1(_04929_),
    .A2(_04942_),
    .A3(_04949_),
    .A4(_04951_),
    .ZN(_04952_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10886_ (.A1(_04666_),
    .A2(_04931_),
    .ZN(_04953_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10887_ (.A1(_04666_),
    .A2(_01990_),
    .B(_04953_),
    .ZN(_04954_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10888_ (.A1(_03857_),
    .A2(_04932_),
    .B1(_04954_),
    .B2(_03697_),
    .C(_02547_),
    .ZN(_04955_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10889_ (.A1(_04952_),
    .A2(_04955_),
    .ZN(_04956_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10890_ (.A1(_03736_),
    .A2(_04932_),
    .ZN(_04957_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10891_ (.A1(\as2650.ivec[3] ),
    .A2(_03736_),
    .B(_04957_),
    .C(_03981_),
    .ZN(_04958_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _10892_ (.A1(_04928_),
    .A2(_04956_),
    .A3(_04958_),
    .ZN(_04959_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10893_ (.A1(_02185_),
    .A2(_04701_),
    .B(_04959_),
    .ZN(_04960_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10894_ (.A1(_03986_),
    .A2(_04960_),
    .ZN(_00344_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10895_ (.A1(_02183_),
    .A2(_04930_),
    .ZN(_04961_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10896_ (.A1(_02195_),
    .A2(_04961_),
    .Z(_04962_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10897_ (.A1(_04179_),
    .A2(_04946_),
    .B(_04271_),
    .ZN(_04963_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _10898_ (.A1(\as2650.addr_buff[0] ),
    .A2(_04214_),
    .A3(_00699_),
    .A4(_04945_),
    .ZN(_04964_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10899_ (.A1(_04682_),
    .A2(_04964_),
    .ZN(_04965_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _10900_ (.A1(_04681_),
    .A2(_04962_),
    .B1(_04963_),
    .B2(_04965_),
    .ZN(_04966_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10901_ (.A1(_02195_),
    .A2(_02182_),
    .A3(_04908_),
    .Z(_04967_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10902_ (.A1(_02184_),
    .A2(_04908_),
    .B(_02196_),
    .ZN(_04968_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _10903_ (.I(_04962_),
    .ZN(_04969_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10904_ (.A1(_00887_),
    .A2(_04969_),
    .ZN(_04970_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _10905_ (.A1(_00888_),
    .A2(_04967_),
    .A3(_04968_),
    .B(_04970_),
    .ZN(_04971_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10906_ (.A1(_02196_),
    .A2(_00603_),
    .ZN(_04972_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10907_ (.A1(_03818_),
    .A2(_04234_),
    .B(_04972_),
    .C(_04541_),
    .ZN(_04973_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10908_ (.A1(_04215_),
    .A2(_00742_),
    .ZN(_04974_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10909_ (.A1(_03841_),
    .A2(_00927_),
    .B(_00747_),
    .ZN(_04975_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10910_ (.A1(_03924_),
    .A2(_04962_),
    .B1(_04974_),
    .B2(_04975_),
    .C(_04367_),
    .ZN(_04976_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10911_ (.A1(_04474_),
    .A2(_04971_),
    .B1(_04973_),
    .B2(_04976_),
    .ZN(_04977_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10912_ (.I(_02559_),
    .Z(_04978_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10913_ (.A1(_03905_),
    .A2(_04234_),
    .B(_04972_),
    .C(_03858_),
    .ZN(_04979_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10914_ (.A1(_04978_),
    .A2(_04969_),
    .B(_04979_),
    .ZN(_04980_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _10915_ (.A1(_04714_),
    .A2(_04977_),
    .B1(_04980_),
    .B2(_00719_),
    .C(_03836_),
    .ZN(_04981_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10916_ (.A1(_00741_),
    .A2(_04966_),
    .B(_04981_),
    .ZN(_04982_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _10917_ (.A1(_00861_),
    .A2(_04559_),
    .ZN(_04983_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10918_ (.I(_00775_),
    .Z(_04984_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _10919_ (.A1(_02042_),
    .A2(_03657_),
    .B1(_04969_),
    .B2(_04983_),
    .C(_04984_),
    .ZN(_04985_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10920_ (.A1(\as2650.ivec[4] ),
    .A2(_04854_),
    .B1(_04856_),
    .B2(_04969_),
    .C(_04698_),
    .ZN(_04986_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10921_ (.A1(_04982_),
    .A2(_04985_),
    .B(_04986_),
    .ZN(_04987_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10922_ (.A1(_02197_),
    .A2(_04701_),
    .B(_04987_),
    .ZN(_04988_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10923_ (.A1(_03986_),
    .A2(_04988_),
    .ZN(_00345_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _10924_ (.I(_02202_),
    .ZN(_04989_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _10925_ (.A1(net65),
    .A2(_02182_),
    .A3(_04930_),
    .ZN(_04990_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10926_ (.A1(_04989_),
    .A2(_04990_),
    .Z(_04991_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10927_ (.A1(_02203_),
    .A2(_02941_),
    .ZN(_04992_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10928_ (.A1(_04082_),
    .A2(_04259_),
    .B(_04992_),
    .ZN(_04993_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10929_ (.A1(_04272_),
    .A2(_00742_),
    .ZN(_04994_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10930_ (.A1(_04688_),
    .A2(_04994_),
    .B(_00747_),
    .ZN(_04995_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _10931_ (.A1(_03925_),
    .A2(_04991_),
    .B1(_04993_),
    .B2(_04704_),
    .C(_04995_),
    .ZN(_04996_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _10932_ (.I(_04991_),
    .Z(_04997_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _10933_ (.A1(_04989_),
    .A2(_04967_),
    .Z(_04998_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10934_ (.A1(_04716_),
    .A2(_04998_),
    .ZN(_04999_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _10935_ (.A1(_00462_),
    .A2(_04997_),
    .B(_04999_),
    .C(_04718_),
    .ZN(_05000_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _10936_ (.A1(_03833_),
    .A2(_04996_),
    .B(_05000_),
    .ZN(_05001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10937_ (.A1(_04250_),
    .A2(_04964_),
    .ZN(_05002_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10938_ (.A1(_04250_),
    .A2(_04964_),
    .ZN(_05003_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10939_ (.A1(_04549_),
    .A2(_05003_),
    .ZN(_05004_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10940_ (.A1(_04632_),
    .A2(_04991_),
    .B1(_05002_),
    .B2(_05004_),
    .ZN(_05005_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10941_ (.A1(_00584_),
    .A2(_04993_),
    .ZN(_05006_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10942_ (.A1(_04978_),
    .A2(_04997_),
    .B(_00542_),
    .ZN(_05007_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _10943_ (.A1(_00514_),
    .A2(_05005_),
    .B1(_05006_),
    .B2(_05007_),
    .C(_03836_),
    .ZN(_05008_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10944_ (.A1(_04616_),
    .A2(_05001_),
    .B(_05008_),
    .ZN(_05009_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _10945_ (.A1(_02065_),
    .A2(_03657_),
    .B1(_04983_),
    .B2(_04997_),
    .C(_04984_),
    .ZN(_05010_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10946_ (.A1(\as2650.ivec[5] ),
    .A2(_04854_),
    .B1(_04856_),
    .B2(_04997_),
    .C(_04698_),
    .ZN(_05011_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10947_ (.A1(_05009_),
    .A2(_05010_),
    .B(_05011_),
    .ZN(_05012_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10948_ (.A1(_02204_),
    .A2(_04701_),
    .B(_05012_),
    .ZN(_05013_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10949_ (.A1(_03986_),
    .A2(_05013_),
    .ZN(_00346_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _10950_ (.A1(_04989_),
    .A2(_04990_),
    .ZN(_05014_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _10951_ (.A1(_02208_),
    .A2(_05014_),
    .Z(_05015_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _10952_ (.I(_05015_),
    .ZN(_05016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10953_ (.A1(_02209_),
    .A2(_00850_),
    .ZN(_05017_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10954_ (.A1(_04082_),
    .A2(_04305_),
    .B(_05017_),
    .ZN(_05018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10955_ (.A1(_04978_),
    .A2(_05018_),
    .ZN(_05019_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10956_ (.A1(_03663_),
    .A2(_05016_),
    .B(_05019_),
    .C(_04244_),
    .ZN(_05020_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10957_ (.A1(_04365_),
    .A2(_05020_),
    .ZN(_05021_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10958_ (.A1(net67),
    .A2(_02202_),
    .A3(_04967_),
    .Z(_05022_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10959_ (.A1(_02203_),
    .A2(_04967_),
    .B(_02209_),
    .ZN(_05023_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _10960_ (.A1(_05022_),
    .A2(_05023_),
    .Z(_05024_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10961_ (.I0(_05016_),
    .I1(_05024_),
    .S(_00461_),
    .Z(_05025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10962_ (.A1(_04704_),
    .A2(_05018_),
    .ZN(_05026_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10963_ (.A1(_04711_),
    .A2(_04049_),
    .B(_04731_),
    .ZN(_05027_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10964_ (.A1(_04245_),
    .A2(_05015_),
    .B1(_05027_),
    .B2(_04400_),
    .C(_03832_),
    .ZN(_05028_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10965_ (.A1(_04368_),
    .A2(_05025_),
    .B1(_05026_),
    .B2(_05028_),
    .ZN(_05029_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _10966_ (.A1(_04249_),
    .A2(_04711_),
    .A3(_04964_),
    .ZN(_05030_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10967_ (.A1(_04289_),
    .A2(_05003_),
    .B(_04863_),
    .ZN(_05031_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _10968_ (.A1(_04681_),
    .A2(_05016_),
    .B1(_05030_),
    .B2(_05031_),
    .C(_00830_),
    .ZN(_05032_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _10969_ (.A1(_00514_),
    .A2(_05029_),
    .B1(_05032_),
    .B2(_04714_),
    .ZN(_05033_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10970_ (.A1(_04595_),
    .A2(_05015_),
    .ZN(_05034_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10971_ (.A1(_04667_),
    .A2(_02095_),
    .B(_04529_),
    .ZN(_05035_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _10972_ (.A1(_05021_),
    .A2(_05033_),
    .B1(_05034_),
    .B2(_05035_),
    .C(_03681_),
    .ZN(_05036_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10973_ (.A1(_03915_),
    .A2(_05016_),
    .B(_04033_),
    .ZN(_05037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _10974_ (.A1(\as2650.ivec[6] ),
    .A2(_04855_),
    .B1(_04857_),
    .B2(_05015_),
    .ZN(_05038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10975_ (.A1(_04523_),
    .A2(_05038_),
    .ZN(_05039_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10976_ (.A1(_05036_),
    .A2(_05037_),
    .B(_05039_),
    .ZN(_05040_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10977_ (.A1(_02210_),
    .A2(_04928_),
    .B(_04702_),
    .ZN(_05041_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10978_ (.A1(_05040_),
    .A2(_05041_),
    .ZN(_00347_));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 _10979_ (.I(_03702_),
    .Z(_05042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _10980_ (.A1(_02208_),
    .A2(_05014_),
    .ZN(_05043_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _10981_ (.A1(_02215_),
    .A2(_05043_),
    .ZN(_05044_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _10982_ (.I(_05044_),
    .Z(_05045_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10983_ (.I0(_02216_),
    .I1(_04336_),
    .S(_03755_),
    .Z(_05046_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _10984_ (.I0(_05045_),
    .I1(_05046_),
    .S(_04978_),
    .Z(_05047_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10985_ (.A1(_04438_),
    .A2(_05030_),
    .B(_04252_),
    .ZN(_05048_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10986_ (.A1(_04438_),
    .A2(_05030_),
    .B(_05048_),
    .ZN(_05049_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10987_ (.A1(_04632_),
    .A2(_05045_),
    .B(_04553_),
    .ZN(_05050_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _10988_ (.A1(_02216_),
    .A2(_05022_),
    .ZN(_05051_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _10989_ (.A1(_02215_),
    .A2(_05022_),
    .Z(_05052_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _10990_ (.A1(_05051_),
    .A2(_05052_),
    .B(_04626_),
    .ZN(_05053_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _10991_ (.A1(_04623_),
    .A2(_05044_),
    .B(_05053_),
    .C(_04640_),
    .ZN(_05054_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _10992_ (.A1(\as2650.addr_buff[4] ),
    .A2(_00723_),
    .B(_00858_),
    .ZN(_05055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _10993_ (.A1(_04774_),
    .A2(_05055_),
    .B(_04885_),
    .ZN(_05056_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _10994_ (.A1(_04126_),
    .A2(_05044_),
    .B1(_05046_),
    .B2(_00859_),
    .C(_05056_),
    .ZN(_05057_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _10995_ (.A1(_00513_),
    .A2(_05054_),
    .A3(_05057_),
    .Z(_05058_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _10996_ (.A1(_05049_),
    .A2(_05050_),
    .B(_05058_),
    .C(_04403_),
    .ZN(_05059_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _10997_ (.A1(_00543_),
    .A2(_05047_),
    .B(_05059_),
    .C(_00861_),
    .ZN(_05060_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _10998_ (.A1(_02118_),
    .A2(_03657_),
    .B1(_04983_),
    .B2(_05045_),
    .C(_00776_),
    .ZN(_05061_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _10999_ (.A1(\as2650.ivec[7] ),
    .A2(_04854_),
    .B1(_04856_),
    .B2(_05045_),
    .C(_04698_),
    .ZN(_05062_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11000_ (.A1(_05060_),
    .A2(_05061_),
    .B(_05062_),
    .ZN(_05063_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11001_ (.A1(_02217_),
    .A2(_04928_),
    .B(_05063_),
    .ZN(_05064_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11002_ (.A1(_05042_),
    .A2(_05064_),
    .ZN(_00348_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _11003_ (.I(net69),
    .ZN(_05065_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _11004_ (.A1(_02215_),
    .A2(_02208_),
    .A3(_05014_),
    .ZN(_05066_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11005_ (.A1(_05065_),
    .A2(_05066_),
    .Z(_05067_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11006_ (.A1(_02224_),
    .A2(_05066_),
    .Z(_05068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11007_ (.A1(_04559_),
    .A2(_05068_),
    .ZN(_05069_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11008_ (.A1(_04667_),
    .A2(_02144_),
    .B(_05069_),
    .C(_04826_),
    .ZN(_05070_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _11009_ (.A1(_04440_),
    .A2(_04076_),
    .B1(_05030_),
    .B2(_04438_),
    .C(_04252_),
    .ZN(_05071_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11010_ (.A1(_04863_),
    .A2(_05067_),
    .B(_00740_),
    .ZN(_05072_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11011_ (.A1(_02224_),
    .A2(_05052_),
    .ZN(_05073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11012_ (.A1(net69),
    .A2(_05052_),
    .ZN(_05074_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11013_ (.A1(_04622_),
    .A2(_05074_),
    .ZN(_05075_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _11014_ (.A1(_04623_),
    .A2(_05068_),
    .B1(_05073_),
    .B2(_05075_),
    .C(_04640_),
    .ZN(_05076_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11015_ (.A1(_02224_),
    .A2(_03817_),
    .ZN(_05077_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11016_ (.A1(_00746_),
    .A2(_00787_),
    .ZN(_05078_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11017_ (.A1(_04440_),
    .A2(_05078_),
    .B(_00535_),
    .ZN(_05079_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _11018_ (.A1(_04126_),
    .A2(_05068_),
    .B1(_05077_),
    .B2(_00859_),
    .C(_05079_),
    .ZN(_05080_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11019_ (.A1(_04553_),
    .A2(_05076_),
    .A3(_05080_),
    .ZN(_05081_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11020_ (.A1(_05071_),
    .A2(_05072_),
    .B(_05081_),
    .C(_04125_),
    .ZN(_05082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11021_ (.A1(_04530_),
    .A2(_05067_),
    .ZN(_05083_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11022_ (.A1(_04669_),
    .A2(_05077_),
    .B(_05083_),
    .C(_04403_),
    .ZN(_05084_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11023_ (.A1(_00834_),
    .A2(_05082_),
    .A3(_05084_),
    .ZN(_05085_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11024_ (.A1(_05070_),
    .A2(_05085_),
    .ZN(_05086_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _11025_ (.A1(_04591_),
    .A2(_05067_),
    .B1(_05086_),
    .B2(_04528_),
    .C(_04592_),
    .ZN(_05087_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _11026_ (.I(_03688_),
    .Z(_05088_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11027_ (.A1(_05065_),
    .A2(_04526_),
    .B(_05087_),
    .C(_05088_),
    .ZN(_00349_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11028_ (.A1(_05065_),
    .A2(_05066_),
    .ZN(_05089_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11029_ (.A1(net71),
    .A2(_05089_),
    .Z(_05090_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11030_ (.I(_05090_),
    .Z(_05091_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11031_ (.A1(_04595_),
    .A2(_05091_),
    .ZN(_05092_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11032_ (.A1(_04667_),
    .A2(_02164_),
    .B(_04529_),
    .ZN(_05093_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11033_ (.A1(_04622_),
    .A2(_05089_),
    .B(_05075_),
    .ZN(_05094_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11034_ (.A1(_02231_),
    .A2(_05094_),
    .Z(_05095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11035_ (.A1(_04245_),
    .A2(_05090_),
    .ZN(_05096_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11036_ (.A1(_02231_),
    .A2(_04024_),
    .Z(_05097_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _11037_ (.A1(_04443_),
    .A2(_05078_),
    .B1(_05097_),
    .B2(_04541_),
    .C(_04367_),
    .ZN(_05098_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11038_ (.A1(_04474_),
    .A2(_05095_),
    .B1(_05096_),
    .B2(_05098_),
    .C(_00740_),
    .ZN(_05099_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11039_ (.A1(_04863_),
    .A2(_05091_),
    .ZN(_05100_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11040_ (.A1(_04682_),
    .A2(_04882_),
    .B(_05100_),
    .C(_04828_),
    .ZN(_05101_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _11041_ (.A1(_00543_),
    .A2(_05099_),
    .A3(_05101_),
    .ZN(_05102_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11042_ (.I0(_05091_),
    .I1(_05097_),
    .S(_03662_),
    .Z(_05103_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11043_ (.A1(_00854_),
    .A2(_05103_),
    .B(_03912_),
    .ZN(_05104_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11044_ (.A1(_05092_),
    .A2(_05093_),
    .B1(_05102_),
    .B2(_05104_),
    .ZN(_05105_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _11045_ (.A1(_04647_),
    .A2(_05091_),
    .B1(_05105_),
    .B2(_04697_),
    .C(_04699_),
    .ZN(_05106_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11046_ (.A1(_02231_),
    .A2(_04928_),
    .B(_04702_),
    .ZN(_05107_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11047_ (.A1(_05106_),
    .A2(_05107_),
    .ZN(_00350_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11048_ (.A1(_00475_),
    .A2(_00895_),
    .B(_00630_),
    .ZN(_05108_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11049_ (.A1(_00769_),
    .A2(_01037_),
    .B(_01031_),
    .C(_00615_),
    .ZN(_05109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11050_ (.A1(_00638_),
    .A2(_00917_),
    .ZN(_05110_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11051_ (.A1(_04416_),
    .A2(_05108_),
    .B1(_05109_),
    .B2(_05110_),
    .ZN(_05111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11052_ (.A1(_03914_),
    .A2(_05111_),
    .ZN(_05112_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11053_ (.A1(_01118_),
    .A2(_02559_),
    .B(_03835_),
    .ZN(_05113_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11054_ (.A1(_00995_),
    .A2(_02522_),
    .B1(_02761_),
    .B2(_02901_),
    .C(_00471_),
    .ZN(_05114_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11055_ (.A1(_00902_),
    .A2(_05113_),
    .B(_05114_),
    .ZN(_05115_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11056_ (.A1(_00884_),
    .A2(_03671_),
    .B(_05115_),
    .ZN(_05116_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11057_ (.A1(_05112_),
    .A2(_05116_),
    .B(_04495_),
    .ZN(_05117_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11058_ (.A1(_00552_),
    .A2(_04421_),
    .B(_03091_),
    .ZN(_05118_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _11059_ (.A1(_00675_),
    .A2(_01013_),
    .A3(_03675_),
    .ZN(_05119_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11060_ (.A1(_02769_),
    .A2(_05118_),
    .A3(_05119_),
    .ZN(_05120_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11061_ (.A1(_02739_),
    .A2(_00503_),
    .A3(_00893_),
    .ZN(_05121_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11062_ (.A1(_03652_),
    .A2(_03713_),
    .Z(_05122_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _11063_ (.A1(_00534_),
    .A2(_00893_),
    .A3(_00982_),
    .ZN(_05123_));
 gf180mcu_fd_sc_mcu7t5v0__oai33_1 _11064_ (.A1(_00523_),
    .A2(_00898_),
    .A3(_05121_),
    .B1(_05122_),
    .B2(_05123_),
    .B3(_00680_),
    .ZN(_05124_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11065_ (.I(net85),
    .ZN(_05125_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11066_ (.A1(\as2650.cycle[9] ),
    .A2(_00902_),
    .A3(_03791_),
    .ZN(_05126_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11067_ (.A1(_00837_),
    .A2(_03723_),
    .ZN(_05127_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11068_ (.A1(_03670_),
    .A2(_05126_),
    .A3(_05127_),
    .ZN(_05128_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11069_ (.A1(_02536_),
    .A2(_05125_),
    .A3(_05128_),
    .ZN(_05129_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _11070_ (.A1(_02765_),
    .A2(_05120_),
    .A3(_05124_),
    .A4(_05129_),
    .Z(_05130_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11071_ (.A1(_05117_),
    .A2(_05130_),
    .Z(_05131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11072_ (.I(_05131_),
    .Z(_05132_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _11073_ (.I(_05132_),
    .Z(_05133_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11074_ (.A1(_04453_),
    .A2(_01094_),
    .ZN(_05134_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11075_ (.I(_00636_),
    .Z(_05135_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11076_ (.I(_00805_),
    .Z(_05136_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11077_ (.A1(_05135_),
    .A2(_01051_),
    .B(_05136_),
    .ZN(_05137_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _11078_ (.A1(_04406_),
    .A2(net82),
    .B1(_05134_),
    .B2(_05137_),
    .C(_03801_),
    .ZN(_05138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _11079_ (.I(_03654_),
    .Z(_05139_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11080_ (.I(_02904_),
    .Z(_05140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11081_ (.I(_00982_),
    .Z(_05141_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11082_ (.I(_05141_),
    .Z(_05142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11083_ (.A1(_00941_),
    .A2(_04585_),
    .ZN(_05143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11084_ (.I(_02530_),
    .Z(_05144_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11085_ (.I(_02530_),
    .Z(_05145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11086_ (.A1(_01760_),
    .A2(_05145_),
    .ZN(_05146_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11087_ (.A1(_01823_),
    .A2(_05144_),
    .B(_01928_),
    .C(_05146_),
    .ZN(_05147_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _11088_ (.A1(_00983_),
    .A2(_05143_),
    .A3(_05147_),
    .ZN(_05148_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11089_ (.I(_00685_),
    .Z(_05149_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _11090_ (.A1(_01146_),
    .A2(_05142_),
    .B(_05148_),
    .C(_05149_),
    .ZN(_05150_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11091_ (.I(_02876_),
    .Z(_05151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11092_ (.I(_00670_),
    .Z(_05152_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11093_ (.A1(_05151_),
    .A2(_01070_),
    .B(_05152_),
    .ZN(_05153_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _11094_ (.A1(_03155_),
    .A2(_05140_),
    .B1(_05150_),
    .B2(_05153_),
    .C(_03654_),
    .ZN(_05154_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _11095_ (.A1(_02857_),
    .A2(_05139_),
    .B(_03666_),
    .C(_05154_),
    .ZN(_05155_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11096_ (.I(_03749_),
    .Z(_05156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11097_ (.A1(_01225_),
    .A2(_05156_),
    .ZN(_05157_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11098_ (.A1(_00914_),
    .A2(_05157_),
    .ZN(_05158_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _11099_ (.A1(_00455_),
    .A2(_04929_),
    .B(_05155_),
    .C(_05158_),
    .ZN(_05159_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11100_ (.A1(_02172_),
    .A2(_01774_),
    .ZN(_05160_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11101_ (.A1(_01777_),
    .A2(_05160_),
    .ZN(_05161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11102_ (.A1(_01822_),
    .A2(_02252_),
    .B(_05161_),
    .ZN(_05162_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11103_ (.I(_05162_),
    .Z(_05163_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11104_ (.A1(_01769_),
    .A2(_01773_),
    .Z(_05164_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11105_ (.I(_05164_),
    .Z(_05165_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _11106_ (.I(_02033_),
    .Z(_05166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11107_ (.A1(\as2650.stack[13][0] ),
    .A2(_05166_),
    .ZN(_05167_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11108_ (.I(_01961_),
    .Z(_05168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11109_ (.I(_02131_),
    .Z(_05169_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11110_ (.I(_02132_),
    .Z(_05170_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _11111_ (.A1(\as2650.stack[14][0] ),
    .A2(_05168_),
    .B1(_05169_),
    .B2(\as2650.stack[15][0] ),
    .C1(\as2650.stack[12][0] ),
    .C2(_05170_),
    .ZN(_05171_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11112_ (.A1(_05165_),
    .A2(_05167_),
    .A3(_05171_),
    .ZN(_05172_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11113_ (.A1(_01808_),
    .A2(_01774_),
    .Z(_05173_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11114_ (.I(_05173_),
    .Z(_05174_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11115_ (.I(_02035_),
    .Z(_05175_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11116_ (.A1(\as2650.stack[11][0] ),
    .A2(_05175_),
    .ZN(_05176_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11117_ (.I(_02137_),
    .Z(_05177_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _11118_ (.A1(\as2650.stack[9][0] ),
    .A2(_05177_),
    .B1(_05170_),
    .B2(\as2650.stack[8][0] ),
    .C1(\as2650.stack[10][0] ),
    .C2(_05168_),
    .ZN(_05178_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11119_ (.A1(_05174_),
    .A2(_05176_),
    .A3(_05178_),
    .ZN(_05179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11120_ (.A1(_05172_),
    .A2(_05179_),
    .ZN(_05180_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11121_ (.I(_02083_),
    .Z(_05181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11122_ (.A1(\as2650.stack[5][0] ),
    .A2(_05181_),
    .ZN(_05182_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _11123_ (.A1(\as2650.stack[6][0] ),
    .A2(_05168_),
    .B1(_02004_),
    .B2(\as2650.stack[7][0] ),
    .C1(\as2650.stack[4][0] ),
    .C2(_02005_),
    .ZN(_05183_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11124_ (.A1(_05165_),
    .A2(_05182_),
    .A3(_05183_),
    .ZN(_05184_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11125_ (.I(_05173_),
    .Z(_05185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11126_ (.I(_02132_),
    .Z(_05186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11127_ (.A1(\as2650.stack[0][0] ),
    .A2(_05186_),
    .ZN(_05187_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11128_ (.A1(\as2650.stack[2][0] ),
    .A2(_05168_),
    .B1(_05169_),
    .B2(\as2650.stack[3][0] ),
    .ZN(_05188_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11129_ (.A1(\as2650.stack[1][0] ),
    .A2(_05177_),
    .ZN(_05189_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _11130_ (.A1(_05185_),
    .A2(_05187_),
    .A3(_05188_),
    .A4(_05189_),
    .ZN(_05190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11131_ (.I(_05162_),
    .Z(_05191_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11132_ (.A1(_05184_),
    .A2(_05190_),
    .B(_05191_),
    .ZN(_05192_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11133_ (.A1(_05163_),
    .A2(_05180_),
    .B(_05192_),
    .ZN(_05193_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11134_ (.I(_04495_),
    .Z(_05194_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11135_ (.I(_05194_),
    .Z(_05195_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _11136_ (.A1(_05138_),
    .A2(_05159_),
    .B1(_05193_),
    .B2(_05195_),
    .C(_05131_),
    .ZN(_05196_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _11137_ (.A1(_01830_),
    .A2(_05133_),
    .B(_05196_),
    .C(_05088_),
    .ZN(_00351_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11138_ (.I(_04420_),
    .Z(_05197_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11139_ (.I(_04063_),
    .Z(_05198_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _11140_ (.A1(_04103_),
    .A2(_01204_),
    .A3(_01205_),
    .ZN(_05199_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _11141_ (.A1(_05198_),
    .A2(_01199_),
    .B(_05199_),
    .C(_04420_),
    .ZN(_05200_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _11142_ (.A1(_05197_),
    .A2(net81),
    .B(_03868_),
    .C(_05200_),
    .ZN(_05201_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11143_ (.I0(_01845_),
    .I1(_01822_),
    .S(_00938_),
    .Z(_05202_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11144_ (.I(_00940_),
    .Z(_05203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11145_ (.A1(_05203_),
    .A2(_04612_),
    .ZN(_05204_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11146_ (.A1(_02741_),
    .A2(_05202_),
    .B(_05204_),
    .C(_02749_),
    .ZN(_05205_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11147_ (.A1(_01237_),
    .A2(_00983_),
    .B(_05205_),
    .C(_00685_),
    .ZN(_05206_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11148_ (.A1(_00830_),
    .A2(_05835_),
    .B(_05206_),
    .ZN(_05207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11149_ (.A1(_02879_),
    .A2(_05207_),
    .ZN(_05208_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11150_ (.A1(_01212_),
    .A2(_00963_),
    .B(_05208_),
    .C(_02888_),
    .ZN(_05209_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11151_ (.A1(_04501_),
    .A2(_02848_),
    .B(_03697_),
    .C(_05209_),
    .ZN(_05210_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _11152_ (.A1(_00454_),
    .A2(_00467_),
    .B1(_03866_),
    .B2(_03155_),
    .C(_05210_),
    .ZN(_05211_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11153_ (.A1(_05201_),
    .A2(_05211_),
    .B(_04447_),
    .ZN(_05212_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11154_ (.I(_05131_),
    .Z(_05213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _11155_ (.I(_05191_),
    .Z(_05214_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11156_ (.I(_05164_),
    .Z(_05215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11157_ (.I(_05215_),
    .Z(_05216_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11158_ (.I(_02008_),
    .Z(_05217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11159_ (.A1(\as2650.stack[13][1] ),
    .A2(_05217_),
    .ZN(_05218_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11160_ (.I(_02087_),
    .Z(_05219_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11161_ (.I(_02089_),
    .Z(_05220_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11162_ (.I(_02090_),
    .Z(_05221_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _11163_ (.A1(\as2650.stack[14][1] ),
    .A2(_05219_),
    .B1(_05220_),
    .B2(\as2650.stack[15][1] ),
    .C1(\as2650.stack[12][1] ),
    .C2(_05221_),
    .ZN(_05222_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11164_ (.A1(_05216_),
    .A2(_05218_),
    .A3(_05222_),
    .ZN(_05223_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11165_ (.I(_05173_),
    .Z(_05224_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11166_ (.I(_02021_),
    .Z(_05225_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11167_ (.A1(\as2650.stack[11][1] ),
    .A2(_05225_),
    .ZN(_05226_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11168_ (.I(_02126_),
    .Z(_05227_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _11169_ (.A1(\as2650.stack[9][1] ),
    .A2(_05227_),
    .B1(_05221_),
    .B2(\as2650.stack[8][1] ),
    .C1(\as2650.stack[10][1] ),
    .C2(_05219_),
    .ZN(_05228_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11170_ (.A1(_05224_),
    .A2(_05226_),
    .A3(_05228_),
    .ZN(_05229_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11171_ (.A1(_05223_),
    .A2(_05229_),
    .ZN(_05230_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11172_ (.I(_02025_),
    .Z(_05231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11173_ (.A1(\as2650.stack[5][1] ),
    .A2(_05231_),
    .ZN(_05232_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11174_ (.I(_02129_),
    .Z(_05233_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11175_ (.I(_02131_),
    .Z(_05234_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _11176_ (.A1(\as2650.stack[6][1] ),
    .A2(_05233_),
    .B1(_05234_),
    .B2(\as2650.stack[7][1] ),
    .C1(\as2650.stack[4][1] ),
    .C2(_05186_),
    .ZN(_05235_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11177_ (.A1(_05216_),
    .A2(_05232_),
    .A3(_05235_),
    .ZN(_05236_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11178_ (.I(_02061_),
    .Z(_05237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11179_ (.A1(\as2650.stack[0][1] ),
    .A2(_05237_),
    .ZN(_05238_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11180_ (.I(_02129_),
    .Z(_05239_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11181_ (.A1(\as2650.stack[2][1] ),
    .A2(_05239_),
    .B1(_05234_),
    .B2(\as2650.stack[3][1] ),
    .ZN(_05240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11182_ (.A1(\as2650.stack[1][1] ),
    .A2(_05166_),
    .ZN(_05241_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _11183_ (.A1(_05185_),
    .A2(_05238_),
    .A3(_05240_),
    .A4(_05241_),
    .ZN(_05242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11184_ (.I(_05162_),
    .Z(_05243_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11185_ (.A1(_05236_),
    .A2(_05242_),
    .B(_05243_),
    .ZN(_05244_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11186_ (.I(_00914_),
    .Z(_05245_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _11187_ (.A1(_05214_),
    .A2(_05230_),
    .B(_05244_),
    .C(_05245_),
    .ZN(_05246_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11188_ (.A1(_05213_),
    .A2(_05246_),
    .ZN(_05247_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11189_ (.I(_00507_),
    .Z(_05248_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _11190_ (.A1(_01851_),
    .A2(_05133_),
    .B1(_05212_),
    .B2(_05247_),
    .C(_05248_),
    .ZN(_00352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11191_ (.A1(_04453_),
    .A2(_01254_),
    .ZN(_05249_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11192_ (.A1(_05198_),
    .A2(_01260_),
    .B(_05249_),
    .C(_05136_),
    .ZN(_05250_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _11193_ (.A1(_00806_),
    .A2(net80),
    .B(_04161_),
    .C(_05250_),
    .ZN(_05251_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11194_ (.I(_00434_),
    .Z(_05252_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11195_ (.I(_02749_),
    .Z(_05253_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11196_ (.I0(_01861_),
    .I1(_01936_),
    .S(_00938_),
    .Z(_05254_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11197_ (.A1(_05203_),
    .A2(_04664_),
    .ZN(_05255_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11198_ (.A1(_02741_),
    .A2(_05254_),
    .B(_05255_),
    .C(_05141_),
    .ZN(_05256_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11199_ (.A1(_01313_),
    .A2(_05253_),
    .B(_05256_),
    .C(_02868_),
    .ZN(_05257_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11200_ (.A1(_03155_),
    .A2(_05149_),
    .B(_05257_),
    .C(_02879_),
    .ZN(_05258_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11201_ (.A1(_05252_),
    .A2(_02879_),
    .B(_05258_),
    .ZN(_05259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11202_ (.A1(_02888_),
    .A2(_05259_),
    .ZN(_05260_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11203_ (.A1(_04503_),
    .A2(_02848_),
    .B(_05260_),
    .ZN(_05261_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11204_ (.I(_00913_),
    .Z(_05262_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11205_ (.A1(_00441_),
    .A2(_00907_),
    .B(_05262_),
    .ZN(_05263_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _11206_ (.A1(_00450_),
    .A2(_03837_),
    .B1(_03810_),
    .B2(_05261_),
    .C(_05263_),
    .ZN(_05264_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11207_ (.I(_05215_),
    .Z(_05265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11208_ (.I(_02394_),
    .Z(_05266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11209_ (.A1(\as2650.stack[13][2] ),
    .A2(_05266_),
    .ZN(_05267_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11210_ (.I(_02059_),
    .Z(_05268_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11211_ (.I(_02061_),
    .Z(_05269_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _11212_ (.A1(\as2650.stack[14][2] ),
    .A2(_05268_),
    .B1(_05175_),
    .B2(\as2650.stack[15][2] ),
    .C1(\as2650.stack[12][2] ),
    .C2(_05269_),
    .ZN(_05270_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11213_ (.A1(_05265_),
    .A2(_05267_),
    .A3(_05270_),
    .ZN(_05271_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11214_ (.I(_05173_),
    .Z(_05272_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11215_ (.I(_02004_),
    .Z(_05273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11216_ (.A1(\as2650.stack[11][2] ),
    .A2(_05273_),
    .ZN(_05274_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11217_ (.I(_02080_),
    .Z(_05275_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11218_ (.I(_02059_),
    .Z(_05276_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _11219_ (.A1(\as2650.stack[9][2] ),
    .A2(_05181_),
    .B1(_05275_),
    .B2(\as2650.stack[8][2] ),
    .C1(\as2650.stack[10][2] ),
    .C2(_05276_),
    .ZN(_05277_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11220_ (.A1(_05272_),
    .A2(_05274_),
    .A3(_05277_),
    .ZN(_05278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11221_ (.A1(_05271_),
    .A2(_05278_),
    .ZN(_05279_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11222_ (.I(_05215_),
    .Z(_05280_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11223_ (.A1(\as2650.stack[5][2] ),
    .A2(_05266_),
    .ZN(_05281_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11224_ (.I(_02082_),
    .Z(_05282_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _11225_ (.A1(\as2650.stack[6][2] ),
    .A2(_05282_),
    .B1(_01815_),
    .B2(\as2650.stack[7][2] ),
    .C1(\as2650.stack[4][2] ),
    .C2(_02254_),
    .ZN(_05283_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11226_ (.A1(_05280_),
    .A2(_05281_),
    .A3(_05283_),
    .ZN(_05284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11227_ (.A1(\as2650.stack[0][2] ),
    .A2(_05237_),
    .ZN(_05285_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11228_ (.I(_02082_),
    .Z(_05286_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11229_ (.I(_01814_),
    .Z(_05287_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11230_ (.A1(\as2650.stack[2][2] ),
    .A2(_05286_),
    .B1(_05287_),
    .B2(\as2650.stack[3][2] ),
    .ZN(_05288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11231_ (.A1(\as2650.stack[1][2] ),
    .A2(_05231_),
    .ZN(_05289_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _11232_ (.A1(_05174_),
    .A2(_05285_),
    .A3(_05288_),
    .A4(_05289_),
    .ZN(_05290_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11233_ (.A1(_05284_),
    .A2(_05290_),
    .B(_05243_),
    .ZN(_05291_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _11234_ (.A1(_05214_),
    .A2(_05279_),
    .B(_05291_),
    .ZN(_05292_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11235_ (.I(_05194_),
    .Z(_05293_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _11236_ (.A1(_05251_),
    .A2(_05264_),
    .B1(_05292_),
    .B2(_05293_),
    .C(_05132_),
    .ZN(_05294_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11237_ (.A1(_05117_),
    .A2(_05130_),
    .ZN(_05295_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11238_ (.I(_00882_),
    .Z(_05296_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11239_ (.A1(_02067_),
    .A2(_05295_),
    .B(_05296_),
    .ZN(_05297_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11240_ (.A1(_05294_),
    .A2(_05297_),
    .ZN(_00353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11241_ (.A1(_04195_),
    .A2(_03958_),
    .ZN(_05298_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11242_ (.A1(_05135_),
    .A2(_01343_),
    .B(_05298_),
    .C(_05136_),
    .ZN(_05299_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _11243_ (.A1(_00806_),
    .A2(_01373_),
    .B(_04161_),
    .C(_05299_),
    .ZN(_05300_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11244_ (.I(_05203_),
    .Z(_05301_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11245_ (.I0(_01872_),
    .I1(_02251_),
    .S(_00939_),
    .Z(_05302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11246_ (.A1(_05301_),
    .A2(_04752_),
    .ZN(_05303_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _11247_ (.A1(_05301_),
    .A2(_05302_),
    .B(_05303_),
    .C(_05253_),
    .ZN(_05304_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11248_ (.A1(_01391_),
    .A2(_05142_),
    .B(_05304_),
    .C(_05149_),
    .ZN(_05305_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11249_ (.A1(_00441_),
    .A2(_05151_),
    .B(_05152_),
    .ZN(_05306_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _11250_ (.A1(_02885_),
    .A2(_02938_),
    .B1(_05305_),
    .B2(_05306_),
    .C(_02902_),
    .ZN(_05307_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _11251_ (.A1(_02865_),
    .A2(_02903_),
    .B(_03666_),
    .C(_05307_),
    .ZN(_05308_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11252_ (.A1(_05252_),
    .A2(_03866_),
    .B(_05262_),
    .ZN(_05309_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _11253_ (.A1(_00452_),
    .A2(_03837_),
    .B(_05308_),
    .C(_05309_),
    .ZN(_05310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11254_ (.A1(\as2650.stack[13][3] ),
    .A2(_05266_),
    .ZN(_05311_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _11255_ (.A1(\as2650.stack[14][3] ),
    .A2(_05268_),
    .B1(_05287_),
    .B2(\as2650.stack[15][3] ),
    .C1(\as2650.stack[12][3] ),
    .C2(_05269_),
    .ZN(_05312_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11256_ (.A1(_05265_),
    .A2(_05311_),
    .A3(_05312_),
    .ZN(_05313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11257_ (.A1(\as2650.stack[11][3] ),
    .A2(_05273_),
    .ZN(_05314_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _11258_ (.A1(\as2650.stack[9][3] ),
    .A2(_05227_),
    .B1(_05275_),
    .B2(\as2650.stack[8][3] ),
    .C1(\as2650.stack[10][3] ),
    .C2(_05268_),
    .ZN(_05315_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11259_ (.A1(_05272_),
    .A2(_05314_),
    .A3(_05315_),
    .ZN(_05316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11260_ (.A1(_05313_),
    .A2(_05316_),
    .ZN(_05317_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11261_ (.A1(\as2650.stack[5][3] ),
    .A2(_05217_),
    .ZN(_05318_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _11262_ (.A1(\as2650.stack[6][3] ),
    .A2(_05282_),
    .B1(_01815_),
    .B2(\as2650.stack[7][3] ),
    .C1(\as2650.stack[4][3] ),
    .C2(_02254_),
    .ZN(_05319_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11263_ (.A1(_05280_),
    .A2(_05318_),
    .A3(_05319_),
    .ZN(_05320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11264_ (.A1(\as2650.stack[0][3] ),
    .A2(_05237_),
    .ZN(_05321_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11265_ (.A1(\as2650.stack[2][3] ),
    .A2(_05286_),
    .B1(_05287_),
    .B2(\as2650.stack[3][3] ),
    .ZN(_05322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11266_ (.A1(\as2650.stack[1][3] ),
    .A2(_05166_),
    .ZN(_05323_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _11267_ (.A1(_05174_),
    .A2(_05321_),
    .A3(_05322_),
    .A4(_05323_),
    .ZN(_05324_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11268_ (.A1(_05320_),
    .A2(_05324_),
    .B(_05243_),
    .ZN(_05325_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11269_ (.A1(_05214_),
    .A2(_05317_),
    .B(_05325_),
    .ZN(_05326_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11270_ (.A1(_05300_),
    .A2(_05310_),
    .B1(_05326_),
    .B2(_05293_),
    .C(_05132_),
    .ZN(_05327_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11271_ (.A1(_02098_),
    .A2(_05295_),
    .B(_05296_),
    .ZN(_05328_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11272_ (.A1(_05327_),
    .A2(_05328_),
    .ZN(_00354_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11273_ (.A1(_05135_),
    .A2(_01413_),
    .ZN(_05329_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11274_ (.A1(_05198_),
    .A2(_01416_),
    .B(_04406_),
    .ZN(_05330_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _11275_ (.A1(_00806_),
    .A2(_01461_),
    .B1(_05329_),
    .B2(_05330_),
    .C(_04161_),
    .ZN(_05331_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11276_ (.A1(net74),
    .A2(_00939_),
    .ZN(_05332_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11277_ (.A1(_01008_),
    .A2(_05145_),
    .ZN(_05333_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11278_ (.A1(_05332_),
    .A2(_05333_),
    .B(_05203_),
    .ZN(_05334_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11279_ (.A1(_00941_),
    .A2(_04801_),
    .B(_05334_),
    .ZN(_05335_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11280_ (.A1(_01724_),
    .A2(_05141_),
    .B(_00685_),
    .ZN(_05336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11281_ (.A1(_05253_),
    .A2(_05335_),
    .B(_05336_),
    .ZN(_05337_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _11282_ (.A1(_05252_),
    .A2(_05151_),
    .B(_05337_),
    .C(_05152_),
    .ZN(_05338_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _11283_ (.A1(_01617_),
    .A2(_02938_),
    .B(_05338_),
    .C(_02902_),
    .ZN(_05339_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _11284_ (.A1(_02850_),
    .A2(_05139_),
    .B(_03666_),
    .C(_05339_),
    .ZN(_05340_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11285_ (.I(_05805_),
    .Z(_05341_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11286_ (.A1(_05341_),
    .A2(_03866_),
    .B(_05262_),
    .ZN(_05342_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _11287_ (.A1(_00437_),
    .A2(_03837_),
    .B(_05340_),
    .C(_05342_),
    .ZN(_05343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11288_ (.A1(\as2650.stack[13][4] ),
    .A2(_05266_),
    .ZN(_05344_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _11289_ (.A1(\as2650.stack[14][4] ),
    .A2(_05286_),
    .B1(_05287_),
    .B2(\as2650.stack[15][4] ),
    .C1(\as2650.stack[12][4] ),
    .C2(_05275_),
    .ZN(_05345_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11290_ (.A1(_05280_),
    .A2(_05344_),
    .A3(_05345_),
    .ZN(_05346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11291_ (.A1(\as2650.stack[11][4] ),
    .A2(_05273_),
    .ZN(_05347_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _11292_ (.A1(\as2650.stack[9][4] ),
    .A2(_05227_),
    .B1(_05275_),
    .B2(\as2650.stack[8][4] ),
    .C1(\as2650.stack[10][4] ),
    .C2(_05268_),
    .ZN(_05348_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11293_ (.A1(_05224_),
    .A2(_05347_),
    .A3(_05348_),
    .ZN(_05349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11294_ (.A1(_05346_),
    .A2(_05349_),
    .ZN(_05350_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11295_ (.A1(\as2650.stack[5][4] ),
    .A2(_05217_),
    .ZN(_05351_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _11296_ (.A1(\as2650.stack[6][4] ),
    .A2(_05282_),
    .B1(_05220_),
    .B2(\as2650.stack[7][4] ),
    .C1(\as2650.stack[4][4] ),
    .C2(_02254_),
    .ZN(_05352_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11297_ (.A1(_05280_),
    .A2(_05351_),
    .A3(_05352_),
    .ZN(_05353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11298_ (.A1(\as2650.stack[0][4] ),
    .A2(_05237_),
    .ZN(_05354_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11299_ (.A1(\as2650.stack[2][4] ),
    .A2(_05286_),
    .B1(_01815_),
    .B2(\as2650.stack[3][4] ),
    .ZN(_05355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11300_ (.A1(\as2650.stack[1][4] ),
    .A2(_05166_),
    .ZN(_05356_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _11301_ (.A1(_05174_),
    .A2(_05354_),
    .A3(_05355_),
    .A4(_05356_),
    .ZN(_05357_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11302_ (.A1(_05353_),
    .A2(_05357_),
    .B(_05243_),
    .ZN(_05358_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11303_ (.A1(_05214_),
    .A2(_05350_),
    .B(_05358_),
    .ZN(_05359_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _11304_ (.A1(_05331_),
    .A2(_05343_),
    .B1(_05359_),
    .B2(_05293_),
    .C(_05132_),
    .ZN(_05360_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11305_ (.A1(_03622_),
    .A2(_05295_),
    .B(_05296_),
    .ZN(_05361_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _11306_ (.A1(_05360_),
    .A2(_05361_),
    .ZN(_00355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11307_ (.A1(_04195_),
    .A2(_01531_),
    .ZN(_05362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11308_ (.A1(_04103_),
    .A2(_01526_),
    .ZN(_05363_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11309_ (.A1(_05362_),
    .A2(_05363_),
    .B(_04420_),
    .ZN(_05364_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11310_ (.A1(_05197_),
    .A2(_01514_),
    .B(_05364_),
    .ZN(_05365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11311_ (.A1(_05341_),
    .A2(_02877_),
    .ZN(_05366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11312_ (.A1(_01894_),
    .A2(_05144_),
    .ZN(_05367_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11313_ (.A1(_02484_),
    .A2(_05144_),
    .B(_05367_),
    .ZN(_05368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11314_ (.A1(_05301_),
    .A2(_04824_),
    .ZN(_05369_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11315_ (.A1(_05301_),
    .A2(_05368_),
    .B(_05369_),
    .C(_05253_),
    .ZN(_05370_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11316_ (.A1(_02223_),
    .A2(_00984_),
    .B(_05370_),
    .C(_05149_),
    .ZN(_05371_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11317_ (.A1(_05366_),
    .A2(_05371_),
    .B(_02938_),
    .ZN(_05372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11318_ (.A1(_01534_),
    .A2(_05140_),
    .ZN(_05373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11319_ (.A1(_02888_),
    .A2(_05373_),
    .ZN(_05374_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _11320_ (.A1(_02554_),
    .A2(_02848_),
    .B1(_05372_),
    .B2(_05374_),
    .C(_03697_),
    .ZN(_05375_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11321_ (.A1(_00428_),
    .A2(_04929_),
    .B1(_05156_),
    .B2(_01422_),
    .ZN(_05376_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11322_ (.A1(_03868_),
    .A2(_05365_),
    .B(_05375_),
    .C(_05376_),
    .ZN(_05377_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11323_ (.A1(_04447_),
    .A2(_05377_),
    .ZN(_05378_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11324_ (.A1(\as2650.stack[13][5] ),
    .A2(_05217_),
    .ZN(_05379_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _11325_ (.A1(\as2650.stack[14][5] ),
    .A2(_05239_),
    .B1(_05220_),
    .B2(\as2650.stack[15][5] ),
    .C1(\as2650.stack[12][5] ),
    .C2(_05221_),
    .ZN(_05380_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11326_ (.A1(_05216_),
    .A2(_05379_),
    .A3(_05380_),
    .ZN(_05381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11327_ (.A1(\as2650.stack[11][5] ),
    .A2(_05225_),
    .ZN(_05382_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _11328_ (.A1(\as2650.stack[9][5] ),
    .A2(_05177_),
    .B1(_05186_),
    .B2(\as2650.stack[8][5] ),
    .C1(\as2650.stack[10][5] ),
    .C2(_05219_),
    .ZN(_05383_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11329_ (.A1(_05224_),
    .A2(_05382_),
    .A3(_05383_),
    .ZN(_05384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11330_ (.A1(_05381_),
    .A2(_05384_),
    .ZN(_05385_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11331_ (.A1(\as2650.stack[5][5] ),
    .A2(_05231_),
    .ZN(_05386_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _11332_ (.A1(\as2650.stack[6][5] ),
    .A2(_05233_),
    .B1(_05169_),
    .B2(\as2650.stack[7][5] ),
    .C1(\as2650.stack[4][5] ),
    .C2(_05170_),
    .ZN(_05387_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11333_ (.A1(_05165_),
    .A2(_05386_),
    .A3(_05387_),
    .ZN(_05388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11334_ (.A1(\as2650.stack[0][5] ),
    .A2(_05269_),
    .ZN(_05389_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11335_ (.A1(\as2650.stack[2][5] ),
    .A2(_05239_),
    .B1(_05234_),
    .B2(\as2650.stack[3][5] ),
    .ZN(_05390_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11336_ (.A1(\as2650.stack[1][5] ),
    .A2(_05181_),
    .ZN(_05391_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _11337_ (.A1(_05185_),
    .A2(_05389_),
    .A3(_05390_),
    .A4(_05391_),
    .ZN(_05392_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11338_ (.A1(_05388_),
    .A2(_05392_),
    .B(_05191_),
    .ZN(_05393_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _11339_ (.A1(_05163_),
    .A2(_05385_),
    .B(_05393_),
    .C(_05245_),
    .ZN(_05394_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11340_ (.A1(_05213_),
    .A2(_05394_),
    .ZN(_05395_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _11341_ (.A1(_01900_),
    .A2(_05133_),
    .B1(_05378_),
    .B2(_05395_),
    .C(_05248_),
    .ZN(_00356_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11342_ (.I(_01606_),
    .ZN(_05396_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11343_ (.A1(_05135_),
    .A2(_01631_),
    .ZN(_05397_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11344_ (.A1(_05198_),
    .A2(_01614_),
    .B(_05197_),
    .ZN(_05398_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _11345_ (.A1(_05197_),
    .A2(_05396_),
    .B1(_05397_),
    .B2(_05398_),
    .ZN(_05399_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11346_ (.A1(net29),
    .A2(_00938_),
    .ZN(_05400_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11347_ (.A1(_05735_),
    .A2(_00939_),
    .B(_05400_),
    .ZN(_05401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11348_ (.A1(_01928_),
    .A2(_05401_),
    .ZN(_05402_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _11349_ (.A1(_01929_),
    .A2(_02847_),
    .B(_05402_),
    .C(_00983_),
    .ZN(_05403_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _11350_ (.A1(_02230_),
    .A2(_05142_),
    .B(_05403_),
    .C(_02868_),
    .ZN(_05404_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11351_ (.A1(_01422_),
    .A2(_05151_),
    .B(_05152_),
    .ZN(_05405_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _11352_ (.A1(_02896_),
    .A2(_05140_),
    .B1(_05404_),
    .B2(_05405_),
    .C(_03654_),
    .ZN(_05406_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _11353_ (.A1(_02854_),
    .A2(_05139_),
    .B(_03653_),
    .C(_05406_),
    .ZN(_05407_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _11354_ (.I(_04495_),
    .Z(_05408_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _11355_ (.A1(_02884_),
    .A2(_05156_),
    .B(_05407_),
    .C(_05408_),
    .ZN(_05409_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_4 _11356_ (.A1(_00424_),
    .A2(_00467_),
    .B1(_03868_),
    .B2(_05399_),
    .C(_05409_),
    .ZN(_05410_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11357_ (.I(_02013_),
    .Z(_05411_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11358_ (.A1(\as2650.stack[13][6] ),
    .A2(_05411_),
    .ZN(_05412_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _11359_ (.A1(\as2650.stack[14][6] ),
    .A2(_05239_),
    .B1(_05220_),
    .B2(\as2650.stack[15][6] ),
    .C1(\as2650.stack[12][6] ),
    .C2(_05221_),
    .ZN(_05413_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11360_ (.A1(_05216_),
    .A2(_05412_),
    .A3(_05413_),
    .ZN(_05414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11361_ (.A1(\as2650.stack[11][6] ),
    .A2(_05225_),
    .ZN(_05415_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _11362_ (.A1(\as2650.stack[9][6] ),
    .A2(_05177_),
    .B1(_05186_),
    .B2(\as2650.stack[8][6] ),
    .C1(\as2650.stack[10][6] ),
    .C2(_05219_),
    .ZN(_05416_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11363_ (.A1(_05224_),
    .A2(_05415_),
    .A3(_05416_),
    .ZN(_05417_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11364_ (.A1(_05414_),
    .A2(_05417_),
    .ZN(_05418_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11365_ (.A1(\as2650.stack[5][6] ),
    .A2(_05231_),
    .ZN(_05419_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _11366_ (.A1(\as2650.stack[6][6] ),
    .A2(_05233_),
    .B1(_05169_),
    .B2(\as2650.stack[7][6] ),
    .C1(\as2650.stack[4][6] ),
    .C2(_05170_),
    .ZN(_05420_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11367_ (.A1(_05165_),
    .A2(_05419_),
    .A3(_05420_),
    .ZN(_05421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11368_ (.A1(\as2650.stack[0][6] ),
    .A2(_05269_),
    .ZN(_05422_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11369_ (.A1(\as2650.stack[2][6] ),
    .A2(_05233_),
    .B1(_05234_),
    .B2(\as2650.stack[3][6] ),
    .ZN(_05423_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11370_ (.A1(\as2650.stack[1][6] ),
    .A2(_05181_),
    .ZN(_05424_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _11371_ (.A1(_05185_),
    .A2(_05422_),
    .A3(_05423_),
    .A4(_05424_),
    .ZN(_05425_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11372_ (.A1(_05421_),
    .A2(_05425_),
    .B(_05191_),
    .ZN(_05426_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _11373_ (.A1(_05163_),
    .A2(_05418_),
    .B(_05426_),
    .C(_05245_),
    .ZN(_05427_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11374_ (.A1(_05213_),
    .A2(_05427_),
    .ZN(_05428_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _11375_ (.A1(_03625_),
    .A2(_05133_),
    .B1(_05410_),
    .B2(_05428_),
    .C(_05248_),
    .ZN(_00357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11376_ (.A1(_04453_),
    .A2(_01702_),
    .ZN(_05429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11377_ (.A1(_04195_),
    .A2(_01713_),
    .ZN(_05430_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11378_ (.A1(_05136_),
    .A2(_05429_),
    .A3(_05430_),
    .ZN(_05431_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11379_ (.A1(_04406_),
    .A2(_03228_),
    .B(_03801_),
    .C(_05431_),
    .ZN(_05432_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11380_ (.A1(_00421_),
    .A2(_04929_),
    .ZN(_05433_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11381_ (.A1(_05727_),
    .A2(_05145_),
    .ZN(_05434_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11382_ (.A1(net77),
    .A2(_05145_),
    .B(_05434_),
    .ZN(_05435_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11383_ (.A1(_02741_),
    .A2(_02966_),
    .ZN(_05436_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11384_ (.A1(_00941_),
    .A2(_05435_),
    .B(_05436_),
    .C(_05141_),
    .ZN(_05437_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11385_ (.A1(_03486_),
    .A2(_05142_),
    .B(_05437_),
    .C(_02868_),
    .ZN(_05438_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11386_ (.A1(_02880_),
    .A2(_05438_),
    .B(_05140_),
    .ZN(_05439_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11387_ (.A1(_02905_),
    .A2(_02883_),
    .B(_05439_),
    .ZN(_05440_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11388_ (.A1(_05139_),
    .A2(_05440_),
    .B(_02943_),
    .ZN(_05441_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _11389_ (.A1(_02784_),
    .A2(_05156_),
    .B1(_03810_),
    .B2(_05441_),
    .C(_05194_),
    .ZN(_05442_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _11390_ (.A1(_05432_),
    .A2(_05433_),
    .A3(_05442_),
    .ZN(_05443_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _11391_ (.A1(_02172_),
    .A2(_02245_),
    .B1(_05160_),
    .B2(_01777_),
    .ZN(_05444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11392_ (.A1(\as2650.stack[3][7] ),
    .A2(_05273_),
    .ZN(_05445_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11393_ (.I(_02016_),
    .Z(_05446_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _11394_ (.A1(\as2650.stack[1][7] ),
    .A2(_05411_),
    .B1(_05446_),
    .B2(\as2650.stack[0][7] ),
    .C1(\as2650.stack[2][7] ),
    .C2(_05276_),
    .ZN(_05447_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11395_ (.A1(_05272_),
    .A2(_05445_),
    .A3(_05447_),
    .ZN(_05448_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11396_ (.A1(\as2650.stack[4][7] ),
    .A2(_05446_),
    .ZN(_05449_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _11397_ (.A1(\as2650.stack[6][7] ),
    .A2(_05276_),
    .B1(_05175_),
    .B2(\as2650.stack[7][7] ),
    .C1(\as2650.stack[5][7] ),
    .C2(_05411_),
    .ZN(_05450_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11398_ (.A1(_05265_),
    .A2(_05449_),
    .A3(_05450_),
    .ZN(_05451_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11399_ (.A1(_05444_),
    .A2(_05448_),
    .A3(_05451_),
    .ZN(_05452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11400_ (.A1(\as2650.stack[14][7] ),
    .A2(_02399_),
    .ZN(_05453_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _11401_ (.A1(\as2650.stack[13][7] ),
    .A2(_05411_),
    .B1(_05446_),
    .B2(\as2650.stack[12][7] ),
    .C1(\as2650.stack[15][7] ),
    .C2(_05225_),
    .ZN(_05454_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11402_ (.A1(_05265_),
    .A2(_05453_),
    .A3(_05454_),
    .ZN(_05455_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11403_ (.A1(\as2650.stack[9][7] ),
    .A2(_03027_),
    .ZN(_05456_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _11404_ (.A1(\as2650.stack[10][7] ),
    .A2(_05276_),
    .B1(_05175_),
    .B2(\as2650.stack[11][7] ),
    .C1(\as2650.stack[8][7] ),
    .C2(_05446_),
    .ZN(_05457_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11405_ (.A1(_05272_),
    .A2(_05456_),
    .A3(_05457_),
    .ZN(_05458_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11406_ (.A1(_05163_),
    .A2(_05455_),
    .A3(_05458_),
    .ZN(_05459_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11407_ (.A1(_02816_),
    .A2(_05452_),
    .A3(_05459_),
    .ZN(_05460_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11408_ (.A1(_05443_),
    .A2(_05460_),
    .B(_05213_),
    .ZN(_05461_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11409_ (.A1(_03285_),
    .A2(_05295_),
    .B(_05296_),
    .ZN(_05462_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11410_ (.A1(_05461_),
    .A2(_05462_),
    .ZN(_00358_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11411_ (.A1(_04412_),
    .A2(_02557_),
    .ZN(_05463_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11412_ (.A1(_02173_),
    .A2(_02857_),
    .B(_03662_),
    .ZN(_05464_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _11413_ (.A1(_01054_),
    .A2(_02561_),
    .A3(_00974_),
    .B1(_05463_),
    .B2(_05464_),
    .ZN(_05465_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11414_ (.A1(_04468_),
    .A2(_00974_),
    .B(_05465_),
    .ZN(_05466_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11415_ (.A1(_02491_),
    .A2(_05466_),
    .B(_05408_),
    .ZN(_05467_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _11416_ (.A1(_00875_),
    .A2(_00855_),
    .A3(_01799_),
    .ZN(_05468_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11417_ (.A1(_04519_),
    .A2(_05468_),
    .B(_00512_),
    .ZN(_05469_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _11418_ (.A1(_03835_),
    .A2(_02740_),
    .B(_02762_),
    .C(_00541_),
    .ZN(_05470_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11419_ (.A1(_04366_),
    .A2(_00788_),
    .B(_02758_),
    .C(_05470_),
    .ZN(_05471_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11420_ (.A1(_02536_),
    .A2(_05471_),
    .ZN(_05472_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11421_ (.A1(_00546_),
    .A2(_01801_),
    .A3(_03729_),
    .ZN(_05473_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _11422_ (.A1(_04048_),
    .A2(_04381_),
    .A3(_05473_),
    .ZN(_05474_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _11423_ (.A1(_02538_),
    .A2(_04380_),
    .A3(_04514_),
    .A4(_05474_),
    .ZN(_05475_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _11424_ (.A1(_02534_),
    .A2(_05469_),
    .A3(_05472_),
    .A4(_05475_),
    .ZN(_05476_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _11425_ (.A1(_02512_),
    .A2(_02528_),
    .A3(_04397_),
    .A4(_05476_),
    .ZN(_05477_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11426_ (.I(_05477_),
    .Z(_05478_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11427_ (.A1(_04033_),
    .A2(_05467_),
    .B(_05478_),
    .ZN(_05479_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11428_ (.A1(_01823_),
    .A2(_05479_),
    .ZN(_05480_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11429_ (.A1(_02491_),
    .A2(_05465_),
    .B(_00840_),
    .ZN(_05481_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11430_ (.A1(_04240_),
    .A2(_05481_),
    .B(_05478_),
    .C(_02173_),
    .ZN(_05482_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11431_ (.A1(_05480_),
    .A2(_05482_),
    .B(_00773_),
    .ZN(_00359_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11432_ (.I(\as2650.r123_2[3][0] ),
    .Z(_05483_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11433_ (.I(_05483_),
    .Z(_00360_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11434_ (.I(\as2650.r123_2[3][1] ),
    .Z(_05484_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11435_ (.I(_05484_),
    .Z(_00361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11436_ (.I(\as2650.r123_2[3][2] ),
    .Z(_05485_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11437_ (.I(_05485_),
    .Z(_00362_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11438_ (.I(\as2650.r123_2[3][3] ),
    .Z(_05486_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11439_ (.I(_05486_),
    .Z(_00363_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11440_ (.I(\as2650.r123_2[3][4] ),
    .Z(_05487_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11441_ (.I(_05487_),
    .Z(_00364_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11442_ (.I(\as2650.r123_2[3][5] ),
    .Z(_05488_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11443_ (.I(_05488_),
    .Z(_00365_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11444_ (.I(\as2650.r123_2[3][6] ),
    .Z(_05489_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11445_ (.I(_05489_),
    .Z(_00366_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11446_ (.I(\as2650.r123_2[3][7] ),
    .Z(_05490_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11447_ (.I(_05490_),
    .Z(_00367_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _11448_ (.A1(_01821_),
    .A2(_01825_),
    .A3(_02246_),
    .ZN(_05491_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11449_ (.I(_05491_),
    .Z(_05492_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11450_ (.I(_05492_),
    .Z(_05493_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11451_ (.I(_05491_),
    .Z(_05494_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11452_ (.A1(\as2650.stack[9][8] ),
    .A2(_05494_),
    .ZN(_05495_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11453_ (.A1(_01767_),
    .A2(_02445_),
    .ZN(_05496_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11454_ (.I(_05496_),
    .Z(_05497_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11455_ (.I(_05497_),
    .Z(_05498_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11456_ (.A1(_02680_),
    .A2(_05493_),
    .B(_05495_),
    .C(_05498_),
    .ZN(_00368_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11457_ (.I(_05491_),
    .Z(_05499_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11458_ (.A1(\as2650.stack[9][9] ),
    .A2(_05499_),
    .ZN(_05500_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11459_ (.A1(_02689_),
    .A2(_05493_),
    .B(_05500_),
    .C(_05498_),
    .ZN(_00369_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11460_ (.A1(\as2650.stack[9][10] ),
    .A2(_05499_),
    .ZN(_05501_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11461_ (.A1(_02692_),
    .A2(_05493_),
    .B(_05501_),
    .C(_05498_),
    .ZN(_00370_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11462_ (.A1(\as2650.stack[9][11] ),
    .A2(_05499_),
    .ZN(_05502_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11463_ (.A1(_02694_),
    .A2(_05493_),
    .B(_05502_),
    .C(_05498_),
    .ZN(_00371_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11464_ (.I(_05492_),
    .Z(_05503_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11465_ (.A1(\as2650.stack[9][12] ),
    .A2(_05499_),
    .ZN(_05504_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11466_ (.I(_05497_),
    .Z(_05505_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11467_ (.A1(_02696_),
    .A2(_05503_),
    .B(_05504_),
    .C(_05505_),
    .ZN(_00372_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11468_ (.A1(\as2650.stack[9][13] ),
    .A2(_05492_),
    .ZN(_05506_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11469_ (.A1(_02700_),
    .A2(_05503_),
    .B(_05506_),
    .C(_05505_),
    .ZN(_00373_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11470_ (.A1(\as2650.stack[9][14] ),
    .A2(_05492_),
    .ZN(_05507_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11471_ (.A1(_02702_),
    .A2(_05503_),
    .B(_05507_),
    .C(_05505_),
    .ZN(_00374_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11472_ (.I(_05496_),
    .Z(_05508_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11473_ (.I(_05508_),
    .Z(_05509_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11474_ (.A1(_02400_),
    .A2(_01816_),
    .A3(_02253_),
    .ZN(_05510_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11475_ (.I(_05510_),
    .Z(_05511_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11476_ (.A1(\as2650.stack[9][0] ),
    .A2(_05511_),
    .ZN(_05512_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _11477_ (.A1(_01840_),
    .A2(_05503_),
    .B(_05505_),
    .ZN(_05513_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11478_ (.A1(_03557_),
    .A2(_05509_),
    .B1(_05512_),
    .B2(_05513_),
    .ZN(_00375_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11479_ (.A1(\as2650.stack[9][1] ),
    .A2(_05511_),
    .ZN(_05514_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11480_ (.I(_05491_),
    .Z(_05515_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11481_ (.I(_05497_),
    .Z(_05516_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11482_ (.A1(_01858_),
    .A2(_05515_),
    .B(_05516_),
    .ZN(_05517_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11483_ (.A1(_03564_),
    .A2(_05509_),
    .B1(_05514_),
    .B2(_05517_),
    .ZN(_00376_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11484_ (.A1(\as2650.stack[9][2] ),
    .A2(_05511_),
    .ZN(_05518_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11485_ (.A1(_01870_),
    .A2(_05515_),
    .B(_05516_),
    .ZN(_05519_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11486_ (.A1(_03569_),
    .A2(_05509_),
    .B1(_05518_),
    .B2(_05519_),
    .ZN(_00377_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11487_ (.A1(\as2650.stack[9][3] ),
    .A2(_05511_),
    .ZN(_05520_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11488_ (.A1(_01881_),
    .A2(_05515_),
    .B(_05516_),
    .ZN(_05521_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11489_ (.A1(_03572_),
    .A2(_05509_),
    .B1(_05520_),
    .B2(_05521_),
    .ZN(_00378_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11490_ (.I(_05497_),
    .Z(_05522_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11491_ (.I(_05510_),
    .Z(_05523_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11492_ (.A1(\as2650.stack[9][4] ),
    .A2(_05523_),
    .ZN(_05524_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11493_ (.A1(_01892_),
    .A2(_05515_),
    .B(_05516_),
    .ZN(_05525_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11494_ (.A1(_03575_),
    .A2(_05522_),
    .B1(_05524_),
    .B2(_05525_),
    .ZN(_00379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11495_ (.A1(\as2650.stack[9][5] ),
    .A2(_05523_),
    .ZN(_05526_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11496_ (.A1(_01906_),
    .A2(_05494_),
    .B(_05508_),
    .ZN(_05527_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11497_ (.A1(_03580_),
    .A2(_05522_),
    .B1(_05526_),
    .B2(_05527_),
    .ZN(_00380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11498_ (.A1(\as2650.stack[9][6] ),
    .A2(_05523_),
    .ZN(_05528_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11499_ (.A1(_01916_),
    .A2(_05494_),
    .B(_05508_),
    .ZN(_05529_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11500_ (.A1(_03583_),
    .A2(_05522_),
    .B1(_05528_),
    .B2(_05529_),
    .ZN(_00381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11501_ (.A1(\as2650.stack[9][7] ),
    .A2(_05523_),
    .ZN(_05530_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11502_ (.A1(_01925_),
    .A2(_05494_),
    .B(_05508_),
    .ZN(_05531_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11503_ (.A1(_03586_),
    .A2(_05522_),
    .B1(_05530_),
    .B2(_05531_),
    .ZN(_00382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11504_ (.A1(_00947_),
    .A2(_01044_),
    .ZN(_05532_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11505_ (.I(_05532_),
    .Z(_05533_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _11506_ (.A1(_00946_),
    .A2(_01044_),
    .B(_01151_),
    .C(_00909_),
    .ZN(_05534_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11507_ (.I(_05534_),
    .Z(_05535_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11508_ (.A1(\as2650.r123[2][0] ),
    .A2(_05535_),
    .ZN(_05536_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _11509_ (.A1(_01403_),
    .A2(_03359_),
    .B1(_05533_),
    .B2(_01141_),
    .C(_05536_),
    .ZN(_00383_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11510_ (.I(_01401_),
    .Z(_05537_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11511_ (.A1(\as2650.r123[2][1] ),
    .A2(_05535_),
    .ZN(_05538_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _11512_ (.A1(_05537_),
    .A2(_03397_),
    .B1(_05533_),
    .B2(_01233_),
    .C(_05538_),
    .ZN(_00384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11513_ (.A1(\as2650.r123[2][2] ),
    .A2(_05535_),
    .ZN(_05539_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _11514_ (.A1(_05537_),
    .A2(_03429_),
    .B1(_05533_),
    .B2(_01305_),
    .C(_05539_),
    .ZN(_00385_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11515_ (.A1(\as2650.r123[2][3] ),
    .A2(_05535_),
    .ZN(_05540_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _11516_ (.A1(_05537_),
    .A2(_03458_),
    .B1(_05533_),
    .B2(_01375_),
    .C(_05540_),
    .ZN(_00386_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11517_ (.I(_05532_),
    .Z(_05541_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11518_ (.I(_05534_),
    .Z(_05542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11519_ (.A1(\as2650.r123[2][4] ),
    .A2(_05542_),
    .ZN(_05543_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _11520_ (.A1(_05537_),
    .A2(_03477_),
    .B1(_05541_),
    .B2(_01462_),
    .C(_05543_),
    .ZN(_00387_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11521_ (.A1(\as2650.r123[2][5] ),
    .A2(_05542_),
    .ZN(_05544_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _11522_ (.A1(_01402_),
    .A2(_03495_),
    .B1(_05541_),
    .B2(_01545_),
    .C(_05544_),
    .ZN(_00388_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11523_ (.A1(\as2650.r123[2][6] ),
    .A2(_05542_),
    .ZN(_05545_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _11524_ (.A1(_01402_),
    .A2(_03502_),
    .B1(_05541_),
    .B2(_01636_),
    .C(_05545_),
    .ZN(_00389_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11525_ (.A1(\as2650.r123[2][7] ),
    .A2(_05542_),
    .ZN(_05546_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _11526_ (.A1(_01402_),
    .A2(_03506_),
    .B1(_05541_),
    .B2(_01718_),
    .C(_05546_),
    .ZN(_00390_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11527_ (.I(net43),
    .ZN(_05547_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11528_ (.A1(_00825_),
    .A2(_01037_),
    .ZN(_05548_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11529_ (.I(_05548_),
    .Z(_05549_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11530_ (.I0(_01225_),
    .I1(_01830_),
    .S(_05549_),
    .Z(_05550_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11531_ (.A1(_00631_),
    .A2(_04417_),
    .B(_04421_),
    .C(_00477_),
    .ZN(_05551_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11532_ (.A1(_00627_),
    .A2(_05551_),
    .ZN(_05552_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _11533_ (.A1(_00607_),
    .A2(_00614_),
    .B(_00884_),
    .C(_00635_),
    .ZN(_05553_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11534_ (.A1(_04348_),
    .A2(_05553_),
    .B(_03671_),
    .ZN(_05554_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _11535_ (.A1(_00876_),
    .A2(_01180_),
    .A3(_03858_),
    .A4(_00501_),
    .ZN(_05555_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _11536_ (.A1(_03676_),
    .A2(_05554_),
    .A3(_05555_),
    .ZN(_05556_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _11537_ (.A1(_03661_),
    .A2(_05552_),
    .A3(_05556_),
    .ZN(_05557_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11538_ (.I(_05557_),
    .Z(_05558_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11539_ (.I0(_05547_),
    .I1(_05550_),
    .S(_05558_),
    .Z(_05559_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11540_ (.A1(_05042_),
    .A2(_05559_),
    .ZN(_00391_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11541_ (.I(net44),
    .ZN(_05560_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11542_ (.I(_05548_),
    .Z(_05561_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11543_ (.I(_05561_),
    .Z(_05562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11544_ (.A1(_01851_),
    .A2(_05562_),
    .ZN(_05563_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11545_ (.A1(_01073_),
    .A2(_05562_),
    .B(_05563_),
    .ZN(_05564_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11546_ (.I0(_05560_),
    .I1(_05564_),
    .S(_05558_),
    .Z(_05565_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11547_ (.A1(_05042_),
    .A2(_05565_),
    .ZN(_00392_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11548_ (.I0(_00441_),
    .I1(_01865_),
    .S(_05549_),
    .Z(_05566_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11549_ (.I0(net45),
    .I1(_05566_),
    .S(_05558_),
    .Z(_05567_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11550_ (.A1(_02570_),
    .A2(_05567_),
    .Z(_05568_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11551_ (.I(_05568_),
    .Z(_00393_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11552_ (.I0(_05252_),
    .I1(_02097_),
    .S(_05561_),
    .Z(_05569_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _11553_ (.I(_05557_),
    .Z(_05570_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11554_ (.I0(net46),
    .I1(_05569_),
    .S(_05570_),
    .Z(_05571_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11555_ (.A1(_02570_),
    .A2(_05571_),
    .Z(_05572_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11556_ (.I(_05572_),
    .Z(_00394_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11557_ (.I0(_05341_),
    .I1(_01421_),
    .S(_05561_),
    .Z(_05573_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11558_ (.I0(net47),
    .I1(_05573_),
    .S(_05570_),
    .Z(_05574_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11559_ (.A1(_02570_),
    .A2(_05574_),
    .Z(_05575_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11560_ (.I(_05575_),
    .Z(_00395_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _11561_ (.I(_00846_),
    .Z(_05576_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11562_ (.A1(_01422_),
    .A2(_05549_),
    .ZN(_05577_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11563_ (.A1(_01900_),
    .A2(_05562_),
    .B(_05577_),
    .ZN(_05578_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11564_ (.I0(net21),
    .I1(_05578_),
    .S(_05570_),
    .Z(_05579_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11565_ (.A1(_05576_),
    .A2(_05579_),
    .Z(_05580_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11566_ (.I(_05580_),
    .Z(_00396_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11567_ (.I(net22),
    .ZN(_05581_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11568_ (.A1(_01911_),
    .A2(_05549_),
    .ZN(_05582_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11569_ (.A1(_01534_),
    .A2(_05562_),
    .B(_05582_),
    .ZN(_05583_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11570_ (.I0(_05581_),
    .I1(_05583_),
    .S(_05558_),
    .Z(_05584_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11571_ (.A1(_05042_),
    .A2(_05584_),
    .ZN(_00397_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11572_ (.I0(_02784_),
    .I1(_03285_),
    .S(_05561_),
    .Z(_05585_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11573_ (.I0(net23),
    .I1(_05585_),
    .S(_05570_),
    .Z(_05586_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11574_ (.A1(_05576_),
    .A2(_05586_),
    .Z(_05587_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11575_ (.I(_05587_),
    .Z(_00398_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11576_ (.I(\as2650.r123[3][0] ),
    .Z(_05588_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11577_ (.I(_05588_),
    .Z(_00399_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11578_ (.I(\as2650.r123[3][1] ),
    .Z(_05589_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11579_ (.I(_05589_),
    .Z(_00400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11580_ (.I(\as2650.r123[3][2] ),
    .Z(_05590_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11581_ (.I(_05590_),
    .Z(_00401_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11582_ (.I(\as2650.r123[3][3] ),
    .Z(_05591_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11583_ (.I(_05591_),
    .Z(_00402_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11584_ (.I(\as2650.r123[3][4] ),
    .Z(_05592_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11585_ (.I(_05592_),
    .Z(_00403_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11586_ (.I(\as2650.r123[3][5] ),
    .Z(_05593_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11587_ (.I(_05593_),
    .Z(_00404_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11588_ (.I(\as2650.r123[3][6] ),
    .Z(_05594_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11589_ (.I(_05594_),
    .Z(_00405_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11590_ (.I(\as2650.r123[3][7] ),
    .Z(_05595_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11591_ (.I(_05595_),
    .Z(_00406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11592_ (.A1(_02850_),
    .A2(_04507_),
    .ZN(_05596_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11593_ (.A1(_03915_),
    .A2(_00802_),
    .B(_05596_),
    .ZN(_00407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11594_ (.A1(_02865_),
    .A2(_04507_),
    .ZN(_05597_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11595_ (.A1(_00877_),
    .A2(_00802_),
    .B(_05597_),
    .ZN(_00408_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _11596_ (.A1(_00838_),
    .A2(_02750_),
    .A3(_02876_),
    .A4(_05144_),
    .ZN(_05598_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11597_ (.A1(_02754_),
    .A2(_02770_),
    .ZN(_05599_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _11598_ (.A1(_00965_),
    .A2(_05122_),
    .A3(_05123_),
    .B(_02776_),
    .ZN(_05600_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _11599_ (.A1(_05598_),
    .A2(_05599_),
    .A3(_05600_),
    .ZN(_05601_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11600_ (.A1(_01368_),
    .A2(_02774_),
    .A3(_03656_),
    .ZN(_05602_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11601_ (.A1(_05121_),
    .A2(_05602_),
    .Z(_05603_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _11602_ (.A1(_02745_),
    .A2(_05119_),
    .A3(_05601_),
    .A4(_05603_),
    .ZN(_05604_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11603_ (.A1(_02746_),
    .A2(_02760_),
    .ZN(_05605_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11604_ (.I(_05605_),
    .ZN(_05606_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _11605_ (.A1(_01117_),
    .A2(_00675_),
    .A3(_02798_),
    .A4(_03675_),
    .ZN(_05607_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _11606_ (.A1(_00959_),
    .A2(_02565_),
    .B1(_04631_),
    .B2(_00552_),
    .C(_02901_),
    .ZN(_05608_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _11607_ (.A1(_02771_),
    .A2(_05606_),
    .A3(_05607_),
    .A4(_05608_),
    .ZN(_05609_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11608_ (.A1(_04640_),
    .A2(_00564_),
    .A3(_02904_),
    .ZN(_05610_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11609_ (.A1(_01063_),
    .A2(_05610_),
    .B(_01065_),
    .ZN(_05611_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _11610_ (.A1(_00919_),
    .A2(_02565_),
    .A3(_01063_),
    .ZN(_05612_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11611_ (.A1(_02763_),
    .A2(_05612_),
    .ZN(_05613_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11612_ (.A1(_02752_),
    .A2(_05613_),
    .ZN(_05614_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _11613_ (.A1(_05604_),
    .A2(_05609_),
    .A3(_05611_),
    .A4(_05614_),
    .ZN(_05615_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11614_ (.A1(_02891_),
    .A2(_04460_),
    .ZN(_05616_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _11615_ (.A1(_05615_),
    .A2(_05616_),
    .ZN(_05617_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11616_ (.A1(_01688_),
    .A2(_01686_),
    .B(_01689_),
    .C(_01505_),
    .ZN(_05618_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _11617_ (.I(_02797_),
    .ZN(_05619_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11618_ (.A1(_01684_),
    .A2(_05619_),
    .B(_01157_),
    .ZN(_05620_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11619_ (.A1(_05618_),
    .A2(_05620_),
    .ZN(_05621_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11620_ (.A1(_03857_),
    .A2(_01346_),
    .A3(_05621_),
    .ZN(_05622_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11621_ (.A1(_01225_),
    .A2(_02905_),
    .ZN(_05623_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11622_ (.A1(_02549_),
    .A2(_02505_),
    .B(_04461_),
    .C(_02869_),
    .ZN(_05624_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11623_ (.A1(_02896_),
    .A2(_02869_),
    .B(_05624_),
    .C(_00963_),
    .ZN(_05625_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _11624_ (.A1(_00628_),
    .A2(_05623_),
    .A3(_05625_),
    .ZN(_05626_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11625_ (.A1(_05622_),
    .A2(_05626_),
    .B(_05408_),
    .ZN(_05627_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _11626_ (.A1(_05293_),
    .A2(_04585_),
    .B(_05627_),
    .C(_05617_),
    .ZN(_05628_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _11627_ (.A1(_01761_),
    .A2(_05617_),
    .B(_05628_),
    .C(_05088_),
    .ZN(_00409_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11628_ (.A1(_01773_),
    .A2(_01965_),
    .ZN(_05629_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11629_ (.A1(_01776_),
    .A2(_05629_),
    .Z(_05630_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11630_ (.A1(_00839_),
    .A2(_03923_),
    .B(_00775_),
    .ZN(_05631_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11631_ (.A1(_01764_),
    .A2(_05164_),
    .ZN(_05632_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11632_ (.A1(_05444_),
    .A2(_05632_),
    .Z(_05633_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11633_ (.A1(_00583_),
    .A2(_02556_),
    .ZN(_05634_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11634_ (.I(_01787_),
    .Z(_05635_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11635_ (.A1(_01324_),
    .A2(_05635_),
    .B(_01929_),
    .C(_04885_),
    .ZN(_05636_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11636_ (.A1(_05635_),
    .A2(_05630_),
    .B(_05636_),
    .ZN(_05637_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11637_ (.A1(_02864_),
    .A2(_05634_),
    .B(_05637_),
    .ZN(_05638_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _11638_ (.A1(_04473_),
    .A2(_00942_),
    .B(_04587_),
    .ZN(_05639_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _11639_ (.I(_02093_),
    .ZN(_05640_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _11640_ (.A1(_02566_),
    .A2(_05638_),
    .B1(_05639_),
    .B2(_05640_),
    .C(_00960_),
    .ZN(_05641_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11641_ (.A1(_05262_),
    .A2(_05633_),
    .B(_05641_),
    .ZN(_05642_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11642_ (.A1(_05630_),
    .A2(_05631_),
    .B1(_05642_),
    .B2(_04984_),
    .ZN(_05643_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11643_ (.A1(_02865_),
    .A2(_01003_),
    .ZN(_05644_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11644_ (.A1(_00969_),
    .A2(_04587_),
    .ZN(_05645_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11645_ (.A1(_05644_),
    .A2(_05645_),
    .ZN(_05646_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11646_ (.A1(_05477_),
    .A2(_05646_),
    .ZN(_05647_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _11647_ (.I0(_05643_),
    .I1(_01785_),
    .S(_05647_),
    .Z(_05648_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11648_ (.A1(_05576_),
    .A2(_05648_),
    .Z(_05649_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11649_ (.I(_05649_),
    .Z(_00410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11650_ (.A1(_00776_),
    .A2(_04559_),
    .ZN(_05650_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _11651_ (.A1(_04503_),
    .A2(_01003_),
    .A3(_05650_),
    .B(_05477_),
    .ZN(_05651_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11652_ (.A1(_02406_),
    .A2(_02298_),
    .ZN(_05652_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11653_ (.A1(_05629_),
    .A2(_05652_),
    .ZN(_05653_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11654_ (.A1(_01764_),
    .A2(_05215_),
    .Z(_05654_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _11655_ (.A1(_01271_),
    .A2(_05635_),
    .B(_01929_),
    .C(_04885_),
    .ZN(_05655_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11656_ (.A1(_05635_),
    .A2(_05653_),
    .B(_05655_),
    .ZN(_05656_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11657_ (.A1(_02860_),
    .A2(_05634_),
    .B(_05656_),
    .ZN(_05657_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _11658_ (.A1(_02003_),
    .A2(_05639_),
    .B1(_05657_),
    .B2(_02566_),
    .C(_00960_),
    .ZN(_05658_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11659_ (.A1(_05245_),
    .A2(_05654_),
    .B(_05658_),
    .ZN(_05659_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11660_ (.A1(_05631_),
    .A2(_05653_),
    .B1(_05659_),
    .B2(_04984_),
    .ZN(_05660_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11661_ (.A1(_05651_),
    .A2(_05660_),
    .ZN(_05661_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11662_ (.A1(_02406_),
    .A2(_05651_),
    .B(_05661_),
    .C(_05088_),
    .ZN(_00411_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11663_ (.A1(_04501_),
    .A2(_01003_),
    .ZN(_05662_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11664_ (.A1(_05645_),
    .A2(_05662_),
    .ZN(_05663_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11665_ (.A1(_05478_),
    .A2(_05663_),
    .ZN(_05664_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _11666_ (.A1(_01981_),
    .A2(_01966_),
    .ZN(_05665_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11667_ (.A1(_02547_),
    .A2(_01798_),
    .ZN(_05666_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _11668_ (.A1(_01209_),
    .A2(_00974_),
    .B1(_00975_),
    .B2(_05665_),
    .C(_00919_),
    .ZN(_05667_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11669_ (.A1(_02557_),
    .A2(_04467_),
    .B(_05667_),
    .ZN(_05668_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_1 _11670_ (.A1(_05282_),
    .A2(_05227_),
    .A3(_05639_),
    .B1(_05668_),
    .B2(_02566_),
    .ZN(_05669_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11671_ (.A1(_02172_),
    .A2(_00839_),
    .B1(_00960_),
    .B2(_05669_),
    .ZN(_05670_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11672_ (.A1(_05665_),
    .A2(_05666_),
    .B1(_05670_),
    .B2(_03981_),
    .ZN(_05671_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _11673_ (.A1(_05478_),
    .A2(_05663_),
    .A3(_05671_),
    .Z(_05672_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11674_ (.A1(_01822_),
    .A2(_05664_),
    .B(_05672_),
    .C(_04757_),
    .ZN(_00412_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _11675_ (.A1(_00537_),
    .A2(_02555_),
    .A3(_00562_),
    .B(_05615_),
    .ZN(_05673_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11676_ (.A1(_02497_),
    .A2(_02550_),
    .B(_04487_),
    .C(_02877_),
    .ZN(_05674_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11677_ (.A1(_05341_),
    .A2(_02877_),
    .B(_05674_),
    .ZN(_05675_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _11678_ (.A1(_02905_),
    .A2(_05675_),
    .B(_05373_),
    .ZN(_05676_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _11679_ (.A1(_02816_),
    .A2(_04824_),
    .B1(_05676_),
    .B2(_02891_),
    .C(_05673_),
    .ZN(_05677_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11680_ (.A1(_01362_),
    .A2(_02791_),
    .Z(_05678_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _11681_ (.A1(_01460_),
    .A2(_05678_),
    .Z(_05679_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11682_ (.A1(_00553_),
    .A2(_05679_),
    .ZN(_05680_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11683_ (.A1(_01895_),
    .A2(_05673_),
    .B1(_05677_),
    .B2(_05680_),
    .C(_05248_),
    .ZN(_00413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11684_ (.A1(_00996_),
    .A2(_02752_),
    .ZN(_05681_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _11685_ (.A1(_04718_),
    .A2(_04503_),
    .A3(_00562_),
    .ZN(_05682_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _11686_ (.A1(_05604_),
    .A2(_05609_),
    .A3(_05681_),
    .A4(_05682_),
    .Z(_05683_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _11687_ (.I(_02505_),
    .Z(_05684_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11688_ (.A1(_01865_),
    .A2(_03833_),
    .B1(_05684_),
    .B2(_04475_),
    .ZN(_05685_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11689_ (.A1(_00562_),
    .A2(_05685_),
    .ZN(_05686_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11690_ (.A1(_05195_),
    .A2(_04664_),
    .B(_05683_),
    .C(_05686_),
    .ZN(_05687_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11691_ (.A1(_01689_),
    .A2(_03228_),
    .ZN(_05688_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _11692_ (.A1(_01688_),
    .A2(_03228_),
    .B(_05688_),
    .C(_00553_),
    .ZN(_05689_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _11693_ (.A1(_01862_),
    .A2(_05683_),
    .B1(_05687_),
    .B2(_05689_),
    .C(_03702_),
    .ZN(_00414_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _11694_ (.A1(_00897_),
    .A2(_00807_),
    .A3(_04558_),
    .A4(_05603_),
    .ZN(_05690_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _11695_ (.A1(_05605_),
    .A2(_05681_),
    .A3(_05690_),
    .ZN(_05691_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _11696_ (.A1(_02745_),
    .A2(_05601_),
    .A3(_05691_),
    .ZN(_05692_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11697_ (.A1(_04447_),
    .A2(_04801_),
    .ZN(_05693_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _11698_ (.A1(_02120_),
    .A2(_00795_),
    .B1(_05684_),
    .B2(_04482_),
    .C(_00840_),
    .ZN(_05694_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _11699_ (.A1(_05194_),
    .A2(_04468_),
    .A3(_02850_),
    .ZN(_05695_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11700_ (.A1(_05695_),
    .A2(_05692_),
    .B(_01230_),
    .ZN(_05696_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _11701_ (.A1(_05692_),
    .A2(_05693_),
    .A3(_05694_),
    .B(_05696_),
    .ZN(_05697_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _11702_ (.A1(_05576_),
    .A2(_05697_),
    .Z(_05698_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _11703_ (.I(_05698_),
    .Z(_00415_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _11704_ (.A1(_05644_),
    .A2(_05692_),
    .Z(_05699_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11705_ (.A1(_02097_),
    .A2(_03833_),
    .B1(_05684_),
    .B2(_04479_),
    .ZN(_05700_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11706_ (.A1(_00840_),
    .A2(_05700_),
    .ZN(_05701_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _11707_ (.A1(_05195_),
    .A2(_04752_),
    .B(_05699_),
    .C(_05701_),
    .ZN(_05702_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _11708_ (.A1(_01873_),
    .A2(_05699_),
    .B(_05702_),
    .C(_04757_),
    .ZN(_00416_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _11709_ (.A1(_05662_),
    .A2(_05692_),
    .Z(_05703_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _11710_ (.A1(_03663_),
    .A2(_04501_),
    .A3(_05684_),
    .ZN(_05704_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11711_ (.A1(_04469_),
    .A2(_05704_),
    .B(_05408_),
    .ZN(_05705_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11712_ (.A1(_05195_),
    .A2(_04612_),
    .B(_05703_),
    .C(_05705_),
    .ZN(_05706_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _11713_ (.A1(_01846_),
    .A2(_05703_),
    .B(_05706_),
    .C(_04757_),
    .ZN(_00417_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11714_ (.A1(_00795_),
    .A2(_04442_),
    .ZN(_05707_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _11715_ (.A1(_03625_),
    .A2(_04489_),
    .B1(_02557_),
    .B2(_04490_),
    .ZN(_05708_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _11716_ (.A1(_02343_),
    .A2(_05707_),
    .A3(_05708_),
    .ZN(_05709_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11717_ (.A1(_02343_),
    .A2(_05707_),
    .B(_02923_),
    .ZN(_05710_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11718_ (.A1(_04702_),
    .A2(_05710_),
    .ZN(_05711_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _11719_ (.A1(_05709_),
    .A2(_05711_),
    .ZN(_00418_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11720_ (.A1(_04489_),
    .A2(_04003_),
    .B(_02343_),
    .ZN(_05712_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _11721_ (.A1(_05725_),
    .A2(_02340_),
    .ZN(_05713_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _11722_ (.A1(_03622_),
    .A2(_00538_),
    .B1(_05713_),
    .B2(_04482_),
    .ZN(_05714_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _11723_ (.A1(net74),
    .A2(_05712_),
    .B(_00846_),
    .ZN(_05715_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _11724_ (.A1(_05712_),
    .A2(_05714_),
    .B(_05715_),
    .ZN(_00419_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11725_ (.D(_00014_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.r123[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11726_ (.D(_00015_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.r123[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11727_ (.D(_00016_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.r123[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11728_ (.D(_00017_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.r123[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11729_ (.D(_00018_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.r123[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11730_ (.D(_00019_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.r123[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11731_ (.D(_00020_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.r123[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11732_ (.D(_00021_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.r123[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11733_ (.D(_00022_),
    .CLK(clknet_leaf_83_wb_clk_i),
    .Q(\as2650.stack[13][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11734_ (.D(_00023_),
    .CLK(clknet_leaf_87_wb_clk_i),
    .Q(\as2650.stack[13][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11735_ (.D(_00024_),
    .CLK(clknet_leaf_87_wb_clk_i),
    .Q(\as2650.stack[13][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11736_ (.D(_00025_),
    .CLK(clknet_leaf_87_wb_clk_i),
    .Q(\as2650.stack[13][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11737_ (.D(_00026_),
    .CLK(clknet_leaf_104_wb_clk_i),
    .Q(\as2650.stack[13][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11738_ (.D(_00027_),
    .CLK(clknet_leaf_104_wb_clk_i),
    .Q(\as2650.stack[13][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11739_ (.D(_00028_),
    .CLK(clknet_leaf_106_wb_clk_i),
    .Q(\as2650.stack[13][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11740_ (.D(_00029_),
    .CLK(clknet_leaf_104_wb_clk_i),
    .Q(\as2650.stack[13][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11741_ (.D(_00030_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.r123[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11742_ (.D(_00031_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.r123[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11743_ (.D(_00032_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.r123[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11744_ (.D(_00033_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.r123[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11745_ (.D(_00034_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.r123[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11746_ (.D(_00035_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.r123[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11747_ (.D(_00036_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.r123[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11748_ (.D(_00037_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.r123[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11749_ (.D(_00038_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.stack[14][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11750_ (.D(_00039_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.stack[14][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11751_ (.D(_00040_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.stack[14][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11752_ (.D(_00041_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.stack[14][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11753_ (.D(_00042_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.stack[14][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11754_ (.D(_00043_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.stack[14][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11755_ (.D(_00044_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.stack[14][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11756_ (.D(_00045_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.stack[13][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11757_ (.D(_00046_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\as2650.stack[13][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11758_ (.D(_00047_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.stack[13][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11759_ (.D(_00048_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.stack[13][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11760_ (.D(_00049_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.stack[13][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11761_ (.D(_00050_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\as2650.stack[13][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11762_ (.D(_00051_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\as2650.stack[13][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11763_ (.D(_00052_),
    .CLK(clknet_leaf_83_wb_clk_i),
    .Q(\as2650.stack[10][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11764_ (.D(_00053_),
    .CLK(clknet_leaf_87_wb_clk_i),
    .Q(\as2650.stack[10][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11765_ (.D(_00054_),
    .CLK(clknet_leaf_87_wb_clk_i),
    .Q(\as2650.stack[10][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11766_ (.D(_00055_),
    .CLK(clknet_leaf_87_wb_clk_i),
    .Q(\as2650.stack[10][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11767_ (.D(_00056_),
    .CLK(clknet_leaf_103_wb_clk_i),
    .Q(\as2650.stack[10][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11768_ (.D(_00057_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.stack[10][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11769_ (.D(_00058_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.stack[10][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11770_ (.D(_00059_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.stack[10][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11771_ (.D(_00060_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.stack[12][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11772_ (.D(_00061_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.stack[12][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11773_ (.D(_00062_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.stack[12][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11774_ (.D(_00063_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.stack[12][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11775_ (.D(_00064_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.stack[12][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11776_ (.D(_00065_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[12][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11777_ (.D(_00066_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.stack[12][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11778_ (.D(_00067_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\as2650.stack[11][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11779_ (.D(_00068_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.stack[11][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11780_ (.D(_00069_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.stack[11][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11781_ (.D(_00070_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.stack[11][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11782_ (.D(_00071_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.stack[11][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11783_ (.D(_00072_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.stack[11][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11784_ (.D(_00073_),
    .CLK(clknet_leaf_11_wb_clk_i),
    .Q(\as2650.stack[11][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11785_ (.D(_00074_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(net77));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11786_ (.D(_00075_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\as2650.stack[14][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11787_ (.D(_00076_),
    .CLK(clknet_leaf_87_wb_clk_i),
    .Q(\as2650.stack[14][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11788_ (.D(_00077_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\as2650.stack[14][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11789_ (.D(_00078_),
    .CLK(clknet_4_11__leaf_wb_clk_i),
    .Q(\as2650.stack[14][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11790_ (.D(_00079_),
    .CLK(clknet_4_9__leaf_wb_clk_i),
    .Q(\as2650.stack[14][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11791_ (.D(_00080_),
    .CLK(clknet_leaf_103_wb_clk_i),
    .Q(\as2650.stack[14][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11792_ (.D(_00081_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.stack[14][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11793_ (.D(_00082_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.stack[14][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11794_ (.D(_00083_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.stack[10][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11795_ (.D(_00084_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.stack[10][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11796_ (.D(_00085_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.stack[10][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11797_ (.D(_00086_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.stack[10][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11798_ (.D(_00087_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.stack[10][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11799_ (.D(_00088_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\as2650.stack[10][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11800_ (.D(_00089_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.stack[10][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11801_ (.D(_00090_),
    .CLK(clknet_leaf_83_wb_clk_i),
    .Q(\as2650.stack[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11802_ (.D(_00091_),
    .CLK(clknet_leaf_86_wb_clk_i),
    .Q(\as2650.stack[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11803_ (.D(_00092_),
    .CLK(clknet_leaf_86_wb_clk_i),
    .Q(\as2650.stack[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11804_ (.D(_00093_),
    .CLK(clknet_leaf_86_wb_clk_i),
    .Q(\as2650.stack[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11805_ (.D(_00094_),
    .CLK(clknet_leaf_105_wb_clk_i),
    .Q(\as2650.stack[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11806_ (.D(_00095_),
    .CLK(clknet_leaf_105_wb_clk_i),
    .Q(\as2650.stack[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11807_ (.D(_00096_),
    .CLK(clknet_leaf_105_wb_clk_i),
    .Q(\as2650.stack[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11808_ (.D(_00097_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\as2650.stack[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11809_ (.D(_00098_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\as2650.stack[0][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11810_ (.D(_00099_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\as2650.stack[0][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11811_ (.D(_00100_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\as2650.stack[0][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11812_ (.D(_00101_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\as2650.stack[0][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11813_ (.D(_00102_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(\as2650.stack[0][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11814_ (.D(_00103_),
    .CLK(clknet_leaf_18_wb_clk_i),
    .Q(\as2650.stack[0][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11815_ (.D(_00104_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\as2650.stack[0][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11816_ (.D(_00105_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\as2650.stack[8][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11817_ (.D(_00106_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.stack[8][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11818_ (.D(_00107_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.stack[8][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11819_ (.D(_00108_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.stack[8][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11820_ (.D(_00109_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\as2650.stack[8][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11821_ (.D(_00110_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\as2650.stack[8][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11822_ (.D(_00111_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\as2650.stack[8][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11823_ (.D(_00112_),
    .CLK(clknet_leaf_112_wb_clk_i),
    .Q(\as2650.stack[7][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11824_ (.D(_00113_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(\as2650.stack[7][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11825_ (.D(_00114_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(\as2650.stack[7][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11826_ (.D(_00115_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\as2650.stack[7][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11827_ (.D(_00116_),
    .CLK(clknet_leaf_112_wb_clk_i),
    .Q(\as2650.stack[7][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11828_ (.D(_00117_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\as2650.stack[7][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11829_ (.D(_00118_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\as2650.stack[7][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11830_ (.D(_00119_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(net75));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11831_ (.D(_00120_),
    .CLK(clknet_leaf_113_wb_clk_i),
    .Q(\as2650.stack[6][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11832_ (.D(_00121_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(\as2650.stack[6][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11833_ (.D(_00122_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(\as2650.stack[6][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11834_ (.D(_00123_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(\as2650.stack[6][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11835_ (.D(_00124_),
    .CLK(clknet_leaf_123_wb_clk_i),
    .Q(\as2650.stack[6][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11836_ (.D(_00125_),
    .CLK(clknet_leaf_113_wb_clk_i),
    .Q(\as2650.stack[6][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11837_ (.D(_00126_),
    .CLK(clknet_leaf_113_wb_clk_i),
    .Q(\as2650.stack[6][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11838_ (.D(_00127_),
    .CLK(clknet_leaf_116_wb_clk_i),
    .Q(\as2650.stack[5][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11839_ (.D(_00128_),
    .CLK(clknet_leaf_114_wb_clk_i),
    .Q(\as2650.stack[5][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11840_ (.D(_00129_),
    .CLK(clknet_leaf_115_wb_clk_i),
    .Q(\as2650.stack[5][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11841_ (.D(_00130_),
    .CLK(clknet_leaf_115_wb_clk_i),
    .Q(\as2650.stack[5][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11842_ (.D(_00131_),
    .CLK(clknet_leaf_114_wb_clk_i),
    .Q(\as2650.stack[5][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11843_ (.D(_00132_),
    .CLK(clknet_leaf_114_wb_clk_i),
    .Q(\as2650.stack[5][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11844_ (.D(_00133_),
    .CLK(clknet_leaf_115_wb_clk_i),
    .Q(\as2650.stack[5][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11845_ (.D(_00134_),
    .CLK(clknet_leaf_109_wb_clk_i),
    .Q(\as2650.stack[4][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11846_ (.D(_00135_),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(\as2650.stack[4][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11847_ (.D(_00136_),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(\as2650.stack[4][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11848_ (.D(_00137_),
    .CLK(clknet_leaf_109_wb_clk_i),
    .Q(\as2650.stack[4][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11849_ (.D(_00138_),
    .CLK(clknet_leaf_111_wb_clk_i),
    .Q(\as2650.stack[4][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11850_ (.D(_00139_),
    .CLK(clknet_4_3__leaf_wb_clk_i),
    .Q(\as2650.stack[4][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11851_ (.D(_00140_),
    .CLK(clknet_leaf_112_wb_clk_i),
    .Q(\as2650.stack[4][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11852_ (.D(_00141_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(\as2650.stack[12][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11853_ (.D(_00142_),
    .CLK(clknet_leaf_82_wb_clk_i),
    .Q(\as2650.stack[12][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11854_ (.D(_00143_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(\as2650.stack[12][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11855_ (.D(_00144_),
    .CLK(clknet_leaf_81_wb_clk_i),
    .Q(\as2650.stack[12][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11856_ (.D(_00145_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\as2650.stack[12][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11857_ (.D(_00146_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.stack[12][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11858_ (.D(_00147_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\as2650.stack[12][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11859_ (.D(_00148_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.stack[12][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11860_ (.D(_00149_),
    .CLK(clknet_leaf_113_wb_clk_i),
    .Q(\as2650.stack[3][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11861_ (.D(_00150_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(\as2650.stack[3][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11862_ (.D(_00151_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(\as2650.stack[3][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11863_ (.D(_00152_),
    .CLK(clknet_leaf_123_wb_clk_i),
    .Q(\as2650.stack[3][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11864_ (.D(_00153_),
    .CLK(clknet_leaf_123_wb_clk_i),
    .Q(\as2650.stack[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11865_ (.D(_00154_),
    .CLK(clknet_leaf_123_wb_clk_i),
    .Q(\as2650.stack[3][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11866_ (.D(_00155_),
    .CLK(clknet_leaf_123_wb_clk_i),
    .Q(\as2650.stack[3][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11867_ (.D(_00156_),
    .CLK(clknet_leaf_126_wb_clk_i),
    .Q(\as2650.stack[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11868_ (.D(_00157_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.stack[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11869_ (.D(_00158_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.stack[2][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11870_ (.D(_00159_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.stack[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11871_ (.D(_00160_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(\as2650.stack[2][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11872_ (.D(_00161_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(\as2650.stack[2][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11873_ (.D(_00162_),
    .CLK(clknet_leaf_125_wb_clk_i),
    .Q(\as2650.stack[2][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11874_ (.D(_00163_),
    .CLK(clknet_leaf_126_wb_clk_i),
    .Q(\as2650.stack[1][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11875_ (.D(_00164_),
    .CLK(clknet_leaf_127_wb_clk_i),
    .Q(\as2650.stack[1][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11876_ (.D(_00165_),
    .CLK(clknet_leaf_127_wb_clk_i),
    .Q(\as2650.stack[1][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11877_ (.D(_00166_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\as2650.stack[1][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11878_ (.D(_00167_),
    .CLK(clknet_leaf_126_wb_clk_i),
    .Q(\as2650.stack[1][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11879_ (.D(_00168_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.stack[1][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11880_ (.D(_00169_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.stack[1][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11881_ (.D(_00170_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\as2650.stack[15][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11882_ (.D(_00171_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.stack[15][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11883_ (.D(_00172_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.stack[15][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11884_ (.D(_00173_),
    .CLK(clknet_leaf_5_wb_clk_i),
    .Q(\as2650.stack[15][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11885_ (.D(_00174_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.stack[15][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11886_ (.D(_00175_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.stack[15][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11887_ (.D(_00176_),
    .CLK(clknet_leaf_127_wb_clk_i),
    .Q(\as2650.stack[15][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11888_ (.D(_00177_),
    .CLK(clknet_4_9__leaf_wb_clk_i),
    .Q(net53));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11889_ (.D(_00178_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(net54));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11890_ (.D(_00179_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\as2650.stack[15][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11891_ (.D(_00180_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.stack[15][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11892_ (.D(_00181_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\as2650.stack[15][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11893_ (.D(_00182_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\as2650.stack[15][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11894_ (.D(_00183_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\as2650.stack[15][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11895_ (.D(_00184_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\as2650.stack[15][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11896_ (.D(_00185_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(\as2650.stack[15][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11897_ (.D(_00186_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(\as2650.stack[15][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11898_ (.D(_00187_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\as2650.stack[8][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11899_ (.D(_00188_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.stack[8][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11900_ (.D(_00189_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.stack[8][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11901_ (.D(_00190_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.stack[8][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11902_ (.D(_00191_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\as2650.stack[8][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11903_ (.D(_00192_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\as2650.stack[8][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11904_ (.D(_00193_),
    .CLK(clknet_leaf_23_wb_clk_i),
    .Q(\as2650.stack[8][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11905_ (.D(_00194_),
    .CLK(clknet_leaf_22_wb_clk_i),
    .Q(\as2650.stack[8][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11906_ (.D(_00195_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\as2650.stack[11][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _11907_ (.D(_00196_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\as2650.stack[11][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11908_ (.D(_00197_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(\as2650.stack[11][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11909_ (.D(_00198_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(\as2650.stack[11][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11910_ (.D(_00199_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(\as2650.stack[11][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11911_ (.D(_00200_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\as2650.stack[11][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11912_ (.D(_00201_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\as2650.stack[11][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11913_ (.D(_00202_),
    .CLK(clknet_leaf_20_wb_clk_i),
    .Q(\as2650.stack[11][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11914_ (.D(_00203_),
    .CLK(clknet_leaf_86_wb_clk_i),
    .Q(\as2650.stack[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11915_ (.D(_00204_),
    .CLK(clknet_leaf_86_wb_clk_i),
    .Q(\as2650.stack[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11916_ (.D(_00205_),
    .CLK(clknet_leaf_84_wb_clk_i),
    .Q(\as2650.stack[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11917_ (.D(_00206_),
    .CLK(clknet_leaf_84_wb_clk_i),
    .Q(\as2650.stack[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11918_ (.D(_00207_),
    .CLK(clknet_leaf_107_wb_clk_i),
    .Q(\as2650.stack[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11919_ (.D(_00208_),
    .CLK(clknet_leaf_106_wb_clk_i),
    .Q(\as2650.stack[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11920_ (.D(_00209_),
    .CLK(clknet_leaf_106_wb_clk_i),
    .Q(\as2650.stack[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11921_ (.D(_00210_),
    .CLK(clknet_leaf_106_wb_clk_i),
    .Q(\as2650.stack[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11922_ (.D(_00211_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.r123_2[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11923_ (.D(_00212_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.r123_2[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11924_ (.D(_00213_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.r123_2[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11925_ (.D(_00214_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.r123_2[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11926_ (.D(_00215_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.r123_2[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11927_ (.D(_00216_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.r123_2[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11928_ (.D(_00217_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.r123_2[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11929_ (.D(_00218_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.r123_2[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11930_ (.D(_00219_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.r123_2[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11931_ (.D(_00220_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.r123_2[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11932_ (.D(_00221_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.r123_2[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11933_ (.D(_00222_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.r123_2[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11934_ (.D(_00223_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.r123_2[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11935_ (.D(_00224_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.r123_2[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11936_ (.D(_00225_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11937_ (.D(_00226_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.r123_2[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11938_ (.D(_00227_),
    .CLK(clknet_leaf_100_wb_clk_i),
    .Q(\as2650.stack[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11939_ (.D(_00228_),
    .CLK(clknet_leaf_98_wb_clk_i),
    .Q(\as2650.stack[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11940_ (.D(_00229_),
    .CLK(clknet_leaf_96_wb_clk_i),
    .Q(\as2650.stack[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11941_ (.D(_00230_),
    .CLK(clknet_leaf_95_wb_clk_i),
    .Q(\as2650.stack[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11942_ (.D(_00231_),
    .CLK(clknet_leaf_94_wb_clk_i),
    .Q(\as2650.stack[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11943_ (.D(_00232_),
    .CLK(clknet_leaf_93_wb_clk_i),
    .Q(\as2650.stack[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11944_ (.D(_00233_),
    .CLK(clknet_leaf_117_wb_clk_i),
    .Q(\as2650.stack[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11945_ (.D(_00234_),
    .CLK(clknet_leaf_117_wb_clk_i),
    .Q(\as2650.stack[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11946_ (.D(_00000_),
    .CLK(clknet_leaf_75_wb_clk_i),
    .Q(\as2650.cycle[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11947_ (.D(_00005_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.cycle[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11948_ (.D(_00006_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.cycle[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11949_ (.D(_00007_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.cycle[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11950_ (.D(_00008_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.cycle[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11951_ (.D(_00009_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.cycle[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11952_ (.D(_00010_),
    .CLK(clknet_4_12__leaf_wb_clk_i),
    .Q(\as2650.cycle[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11953_ (.D(_00011_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.cycle[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _11954_ (.D(_00012_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\as2650.cycle[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11955_ (.D(_00013_),
    .CLK(clknet_leaf_59_wb_clk_i),
    .Q(\as2650.cycle[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11956_ (.D(_00001_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.cycle[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11957_ (.D(_00002_),
    .CLK(clknet_4_13__leaf_wb_clk_i),
    .Q(\as2650.cycle[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11958_ (.D(_00003_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\as2650.cycle[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11959_ (.D(_00004_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.cycle[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11960_ (.D(_00235_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.r123_2[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11961_ (.D(_00236_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.r123_2[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11962_ (.D(_00237_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.r123_2[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11963_ (.D(_00238_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.r123_2[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11964_ (.D(_00239_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.r123_2[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11965_ (.D(_00240_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.r123_2[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11966_ (.D(_00241_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.r123_2[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11967_ (.D(_00242_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.r123_2[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11968_ (.D(_00243_),
    .CLK(clknet_leaf_94_wb_clk_i),
    .Q(\as2650.stack[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11969_ (.D(_00244_),
    .CLK(clknet_leaf_95_wb_clk_i),
    .Q(\as2650.stack[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11970_ (.D(_00245_),
    .CLK(clknet_leaf_96_wb_clk_i),
    .Q(\as2650.stack[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11971_ (.D(_00246_),
    .CLK(clknet_leaf_95_wb_clk_i),
    .Q(\as2650.stack[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11972_ (.D(_00247_),
    .CLK(clknet_leaf_92_wb_clk_i),
    .Q(\as2650.stack[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11973_ (.D(_00248_),
    .CLK(clknet_leaf_93_wb_clk_i),
    .Q(\as2650.stack[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11974_ (.D(_00249_),
    .CLK(clknet_leaf_117_wb_clk_i),
    .Q(\as2650.stack[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11975_ (.D(_00250_),
    .CLK(clknet_leaf_117_wb_clk_i),
    .Q(\as2650.stack[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11976_ (.D(_00251_),
    .CLK(clknet_leaf_94_wb_clk_i),
    .Q(\as2650.stack[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11977_ (.D(_00252_),
    .CLK(clknet_leaf_96_wb_clk_i),
    .Q(\as2650.stack[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11978_ (.D(_00253_),
    .CLK(clknet_leaf_96_wb_clk_i),
    .Q(\as2650.stack[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11979_ (.D(_00254_),
    .CLK(clknet_leaf_95_wb_clk_i),
    .Q(\as2650.stack[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11980_ (.D(_00255_),
    .CLK(clknet_leaf_94_wb_clk_i),
    .Q(\as2650.stack[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11981_ (.D(_00256_),
    .CLK(clknet_leaf_93_wb_clk_i),
    .Q(\as2650.stack[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11982_ (.D(_00257_),
    .CLK(clknet_leaf_118_wb_clk_i),
    .Q(\as2650.stack[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11983_ (.D(_00258_),
    .CLK(clknet_leaf_118_wb_clk_i),
    .Q(\as2650.stack[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11984_ (.D(_00259_),
    .CLK(clknet_leaf_100_wb_clk_i),
    .Q(\as2650.stack[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11985_ (.D(_00260_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\as2650.stack[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11986_ (.D(_00261_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\as2650.stack[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11987_ (.D(_00262_),
    .CLK(clknet_leaf_98_wb_clk_i),
    .Q(\as2650.stack[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11988_ (.D(_00263_),
    .CLK(clknet_leaf_100_wb_clk_i),
    .Q(\as2650.stack[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11989_ (.D(_00264_),
    .CLK(clknet_leaf_102_wb_clk_i),
    .Q(\as2650.stack[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11990_ (.D(_00265_),
    .CLK(clknet_leaf_118_wb_clk_i),
    .Q(\as2650.stack[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11991_ (.D(_00266_),
    .CLK(clknet_leaf_117_wb_clk_i),
    .Q(\as2650.stack[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11992_ (.D(_00267_),
    .CLK(clknet_leaf_98_wb_clk_i),
    .Q(\as2650.stack[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11993_ (.D(_00268_),
    .CLK(clknet_leaf_84_wb_clk_i),
    .Q(\as2650.stack[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11994_ (.D(_00269_),
    .CLK(clknet_leaf_85_wb_clk_i),
    .Q(\as2650.stack[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11995_ (.D(_00270_),
    .CLK(clknet_leaf_84_wb_clk_i),
    .Q(\as2650.stack[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11996_ (.D(_00271_),
    .CLK(clknet_leaf_100_wb_clk_i),
    .Q(\as2650.stack[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11997_ (.D(_00272_),
    .CLK(clknet_leaf_102_wb_clk_i),
    .Q(\as2650.stack[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11998_ (.D(_00273_),
    .CLK(clknet_leaf_107_wb_clk_i),
    .Q(\as2650.stack[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _11999_ (.D(_00274_),
    .CLK(clknet_4_3__leaf_wb_clk_i),
    .Q(\as2650.stack[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12000_ (.D(_00275_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\as2650.ivec[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12001_ (.D(_00276_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(\as2650.ivec[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12002_ (.D(_00277_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(\as2650.ivec[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12003_ (.D(_00278_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(\as2650.ivec[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12004_ (.D(_00279_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\as2650.ivec[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12005_ (.D(_00280_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\as2650.ivec[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12006_ (.D(_00281_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(\as2650.ivec[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12007_ (.D(_00282_),
    .CLK(clknet_leaf_72_wb_clk_i),
    .Q(\as2650.ivec[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12008_ (.D(_00283_),
    .CLK(clknet_leaf_99_wb_clk_i),
    .Q(\as2650.stack[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12009_ (.D(_00284_),
    .CLK(clknet_leaf_85_wb_clk_i),
    .Q(\as2650.stack[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12010_ (.D(_00285_),
    .CLK(clknet_leaf_84_wb_clk_i),
    .Q(\as2650.stack[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12011_ (.D(_00286_),
    .CLK(clknet_leaf_85_wb_clk_i),
    .Q(\as2650.stack[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12012_ (.D(_00287_),
    .CLK(clknet_4_8__leaf_wb_clk_i),
    .Q(\as2650.stack[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12013_ (.D(_00288_),
    .CLK(clknet_leaf_102_wb_clk_i),
    .Q(\as2650.stack[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12014_ (.D(_00289_),
    .CLK(clknet_leaf_107_wb_clk_i),
    .Q(\as2650.stack[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12015_ (.D(_00290_),
    .CLK(clknet_leaf_107_wb_clk_i),
    .Q(\as2650.stack[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12016_ (.D(_00291_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12017_ (.D(_00292_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12018_ (.D(_00293_),
    .CLK(clknet_leaf_58_wb_clk_i),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12019_ (.D(_00294_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12020_ (.D(_00295_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12021_ (.D(_00296_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12022_ (.D(_00297_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12023_ (.D(_00298_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(net34));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12024_ (.D(_00299_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(net35));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12025_ (.D(_00300_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(net36));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12026_ (.D(_00301_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(net37));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12027_ (.D(_00302_),
    .CLK(clknet_leaf_66_wb_clk_i),
    .Q(net38));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12028_ (.D(_00303_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(net39));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12029_ (.D(_00304_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(net40));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12030_ (.D(_00305_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(net41));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12031_ (.D(_00306_),
    .CLK(clknet_leaf_67_wb_clk_i),
    .Q(net42));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12032_ (.D(_00307_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12033_ (.D(_00308_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12034_ (.D(_00309_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\as2650.addr_buff[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12035_ (.D(_00310_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\as2650.addr_buff[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12036_ (.D(_00311_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\as2650.addr_buff[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12037_ (.D(_00312_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\as2650.addr_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12038_ (.D(_00313_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\as2650.addr_buff[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12039_ (.D(_00314_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.addr_buff[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12040_ (.D(_00315_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.addr_buff[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12041_ (.D(_00316_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\as2650.addr_buff[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12042_ (.D(_00317_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\as2650.last_intr ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12043_ (.D(_00318_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\as2650.prefixed ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12044_ (.D(_00319_),
    .CLK(clknet_4_7__leaf_wb_clk_i),
    .Q(\as2650.idx_ctrl[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12045_ (.D(_00320_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.idx_ctrl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12046_ (.D(_00321_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.holding_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12047_ (.D(_00322_),
    .CLK(clknet_4_7__leaf_wb_clk_i),
    .Q(\as2650.holding_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12048_ (.D(_00323_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.holding_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12049_ (.D(_00324_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.holding_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12050_ (.D(_00325_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\as2650.holding_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12051_ (.D(_00326_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.holding_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12052_ (.D(_00327_),
    .CLK(clknet_leaf_79_wb_clk_i),
    .Q(\as2650.holding_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12053_ (.D(_00328_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(\as2650.holding_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12054_ (.D(_00329_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.ins_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12055_ (.D(_00330_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.ins_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12056_ (.D(_00331_),
    .CLK(clknet_leaf_75_wb_clk_i),
    .Q(\as2650.ins_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12057_ (.D(_00332_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.alu_op[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12058_ (.D(_00333_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\as2650.alu_op[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12059_ (.D(_00334_),
    .CLK(clknet_leaf_76_wb_clk_i),
    .Q(\as2650.alu_op[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12060_ (.D(_00335_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(net72));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _12061_ (.D(_00336_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(net55));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _12062_ (.D(_00337_),
    .CLK(clknet_leaf_74_wb_clk_i),
    .Q(net56));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _12063_ (.D(_00338_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(net57));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _12064_ (.D(_00339_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(net58));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _12065_ (.D(_00340_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(net60));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _12066_ (.D(_00341_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(net61));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _12067_ (.D(_00342_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(net62));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12068_ (.D(_00343_),
    .CLK(clknet_leaf_69_wb_clk_i),
    .Q(net63));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _12069_ (.D(_00344_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(net64));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12070_ (.D(_00345_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(net65));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _12071_ (.D(_00346_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(net66));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12072_ (.D(_00347_),
    .CLK(clknet_leaf_70_wb_clk_i),
    .Q(net67));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _12073_ (.D(_00348_),
    .CLK(clknet_leaf_71_wb_clk_i),
    .Q(net68));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _12074_ (.D(_00349_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(net69));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _12075_ (.D(_00350_),
    .CLK(clknet_leaf_68_wb_clk_i),
    .Q(net71));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12076_ (.D(_00351_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.r0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12077_ (.D(_00352_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.r0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12078_ (.D(_00353_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.r0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12079_ (.D(_00354_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.r0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12080_ (.D(_00355_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.r0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12081_ (.D(_00356_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.r0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12082_ (.D(_00357_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\as2650.r0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12083_ (.D(_00358_),
    .CLK(clknet_leaf_26_wb_clk_i),
    .Q(\as2650.r0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12084_ (.D(_00359_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(net48));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12085_ (.D(_00360_),
    .CLK(clknet_leaf_86_wb_clk_i),
    .Q(\as2650.r123_2[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12086_ (.D(_00361_),
    .CLK(clknet_leaf_91_wb_clk_i),
    .Q(\as2650.r123_2[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12087_ (.D(_00362_),
    .CLK(clknet_leaf_120_wb_clk_i),
    .Q(\as2650.r123_2[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12088_ (.D(_00363_),
    .CLK(clknet_leaf_91_wb_clk_i),
    .Q(\as2650.r123_2[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12089_ (.D(_00364_),
    .CLK(clknet_4_0__leaf_wb_clk_i),
    .Q(\as2650.r123_2[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12090_ (.D(_00365_),
    .CLK(clknet_4_2__leaf_wb_clk_i),
    .Q(\as2650.r123_2[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12091_ (.D(_00366_),
    .CLK(clknet_4_2__leaf_wb_clk_i),
    .Q(\as2650.r123_2[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12092_ (.D(_00367_),
    .CLK(clknet_leaf_116_wb_clk_i),
    .Q(\as2650.r123_2[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12093_ (.D(_00368_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\as2650.stack[9][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12094_ (.D(_00369_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.stack[9][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12095_ (.D(_00370_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.stack[9][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12096_ (.D(_00371_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.stack[9][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12097_ (.D(_00372_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.stack[9][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12098_ (.D(_00373_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.stack[9][13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12099_ (.D(_00374_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.stack[9][14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12100_ (.D(_00375_),
    .CLK(clknet_leaf_99_wb_clk_i),
    .Q(\as2650.stack[9][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12101_ (.D(_00376_),
    .CLK(clknet_leaf_97_wb_clk_i),
    .Q(\as2650.stack[9][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12102_ (.D(_00377_),
    .CLK(clknet_leaf_99_wb_clk_i),
    .Q(\as2650.stack[9][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12103_ (.D(_00378_),
    .CLK(clknet_leaf_99_wb_clk_i),
    .Q(\as2650.stack[9][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12104_ (.D(_00379_),
    .CLK(clknet_leaf_102_wb_clk_i),
    .Q(\as2650.stack[9][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12105_ (.D(_00380_),
    .CLK(clknet_leaf_102_wb_clk_i),
    .Q(\as2650.stack[9][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12106_ (.D(_00381_),
    .CLK(clknet_leaf_109_wb_clk_i),
    .Q(\as2650.stack[9][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12107_ (.D(_00382_),
    .CLK(clknet_leaf_109_wb_clk_i),
    .Q(\as2650.stack[9][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12108_ (.D(_00383_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.r123[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12109_ (.D(_00384_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.r123[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12110_ (.D(_00385_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.r123[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12111_ (.D(_00386_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.r123[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12112_ (.D(_00387_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.r123[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12113_ (.D(_00388_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.r123[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12114_ (.D(_00389_),
    .CLK(clknet_4_5__leaf_wb_clk_i),
    .Q(\as2650.r123[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12115_ (.D(_00390_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.r123[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12116_ (.D(_00391_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(net43));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12117_ (.D(_00392_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(net44));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12118_ (.D(_00393_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(net45));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12119_ (.D(_00394_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(net46));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12120_ (.D(_00395_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(net47));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12121_ (.D(_00396_),
    .CLK(clknet_4_12__leaf_wb_clk_i),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12122_ (.D(_00397_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12123_ (.D(_00398_),
    .CLK(clknet_4_12__leaf_wb_clk_i),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12124_ (.D(_00399_),
    .CLK(clknet_leaf_116_wb_clk_i),
    .Q(\as2650.r123[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12125_ (.D(_00400_),
    .CLK(clknet_leaf_119_wb_clk_i),
    .Q(\as2650.r123[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12126_ (.D(_00401_),
    .CLK(clknet_leaf_92_wb_clk_i),
    .Q(\as2650.r123[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12127_ (.D(_00402_),
    .CLK(clknet_leaf_119_wb_clk_i),
    .Q(\as2650.r123[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12128_ (.D(_00403_),
    .CLK(clknet_leaf_120_wb_clk_i),
    .Q(\as2650.r123[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12129_ (.D(_00404_),
    .CLK(clknet_4_10__leaf_wb_clk_i),
    .Q(\as2650.r123[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12130_ (.D(_00405_),
    .CLK(clknet_4_0__leaf_wb_clk_i),
    .Q(\as2650.r123[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12131_ (.D(_00406_),
    .CLK(clknet_leaf_119_wb_clk_i),
    .Q(\as2650.r123[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12132_ (.D(_00407_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\as2650.ins_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _12133_ (.D(_00408_),
    .CLK(clknet_leaf_73_wb_clk_i),
    .Q(\as2650.ins_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _12134_ (.D(_00409_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(net78));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _12135_ (.D(_00410_),
    .CLK(clknet_leaf_79_wb_clk_i),
    .Q(net73));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _12136_ (.D(_00411_),
    .CLK(clknet_leaf_79_wb_clk_i),
    .Q(net70));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _12137_ (.D(_00412_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(net59));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _12138_ (.D(_00413_),
    .CLK(clknet_4_9__leaf_wb_clk_i),
    .Q(net52));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _12139_ (.D(_00414_),
    .CLK(clknet_leaf_78_wb_clk_i),
    .Q(net49));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _12140_ (.D(_00415_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(net51));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _12141_ (.D(_00416_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(net50));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _12142_ (.D(_00417_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(net79));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _12143_ (.D(_00418_),
    .CLK(clknet_leaf_77_wb_clk_i),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffq_4 _12144_ (.D(_00419_),
    .CLK(clknet_leaf_79_wb_clk_i),
    .Q(net74));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12218_ (.I(net86),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12219_ (.I(net86),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12220_ (.I(net86),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12221_ (.I(net86),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12222_ (.I(net87),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12223_ (.I(net88),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12224_ (.I(net88),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _12225_ (.I(net29),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_wb_clk_i (.I(wb_clk_i),
    .Z(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_0_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_1_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_2_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_3_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_4_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_5_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_6_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_7_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_0__f_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_4_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_10__f_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_4_10__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_11__f_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_4_11__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_12__f_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_4_12__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_13__f_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_4_13__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_14__f_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_4_14__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_15__f_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_4_15__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_1__f_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_4_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_2__f_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_4_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_3__f_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_4_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_4__f_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_4_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_5__f_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_4_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_6__f_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_4_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_7__f_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_4_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_8__f_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_4_8__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_4_9__f_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_4_9__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_0_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_100_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_100_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_102_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_102_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_103_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_103_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_104_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_104_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_105_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_105_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_106_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_106_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_107_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_107_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_109_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_109_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_10_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_10_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_111_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_111_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_112_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_112_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_113_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_113_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_114_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_114_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_115_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_115_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_116_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_116_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_117_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_117_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_118_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_118_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_119_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_119_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_11_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_11_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_120_wb_clk_i (.I(clknet_4_2__leaf_wb_clk_i),
    .Z(clknet_leaf_120_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_123_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_123_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_125_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_125_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_126_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_126_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_127_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_127_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_12_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_12_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_13_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_13_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_14_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_14_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_15_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_16_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_16_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_17_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_17_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_18_wb_clk_i (.I(clknet_4_0__leaf_wb_clk_i),
    .Z(clknet_leaf_18_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_19_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_19_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_1_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_20_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_20_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_21_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_21_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_22_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_22_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_23_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_23_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_24_wb_clk_i (.I(clknet_4_3__leaf_wb_clk_i),
    .Z(clknet_leaf_24_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_25_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_26_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_26_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_27_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_28_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_28_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_29_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_29_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_2_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_31_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_32_wb_clk_i (.I(clknet_4_6__leaf_wb_clk_i),
    .Z(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_33_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_34_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_35_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_35_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_36_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_37_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_38_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_39_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_3_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_40_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_41_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_42_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_43_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_44_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_46_wb_clk_i (.I(clknet_4_5__leaf_wb_clk_i),
    .Z(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_48_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_49_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_4_wb_clk_i (.I(clknet_4_1__leaf_wb_clk_i),
    .Z(clknet_leaf_4_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_50_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_52_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_53_wb_clk_i (.I(clknet_4_7__leaf_wb_clk_i),
    .Z(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_58_wb_clk_i (.I(clknet_4_13__leaf_wb_clk_i),
    .Z(clknet_leaf_58_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_59_wb_clk_i (.I(clknet_4_12__leaf_wb_clk_i),
    .Z(clknet_leaf_59_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_5_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_5_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_60_wb_clk_i (.I(clknet_4_13__leaf_wb_clk_i),
    .Z(clknet_leaf_60_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_61_wb_clk_i (.I(clknet_4_13__leaf_wb_clk_i),
    .Z(clknet_leaf_61_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_63_wb_clk_i (.I(clknet_4_13__leaf_wb_clk_i),
    .Z(clknet_leaf_63_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_64_wb_clk_i (.I(clknet_4_13__leaf_wb_clk_i),
    .Z(clknet_leaf_64_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_65_wb_clk_i (.I(clknet_4_15__leaf_wb_clk_i),
    .Z(clknet_leaf_65_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_66_wb_clk_i (.I(clknet_4_15__leaf_wb_clk_i),
    .Z(clknet_leaf_66_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_67_wb_clk_i (.I(clknet_4_15__leaf_wb_clk_i),
    .Z(clknet_leaf_67_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_68_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_68_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_69_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_69_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_6_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_6_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_70_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_70_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_71_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_71_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_72_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_72_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_73_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_73_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_74_wb_clk_i (.I(clknet_4_15__leaf_wb_clk_i),
    .Z(clknet_leaf_74_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_75_wb_clk_i (.I(clknet_4_14__leaf_wb_clk_i),
    .Z(clknet_leaf_75_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_76_wb_clk_i (.I(clknet_4_12__leaf_wb_clk_i),
    .Z(clknet_leaf_76_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_77_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_77_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_78_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_78_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_79_wb_clk_i (.I(clknet_4_9__leaf_wb_clk_i),
    .Z(clknet_leaf_79_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_7_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_7_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_81_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_81_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_82_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_82_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_83_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_83_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_84_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_84_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_85_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_85_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_86_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_86_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_87_wb_clk_i (.I(clknet_4_11__leaf_wb_clk_i),
    .Z(clknet_leaf_87_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_8_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_8_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_91_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_91_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_92_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_92_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_93_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_93_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_94_wb_clk_i (.I(clknet_4_8__leaf_wb_clk_i),
    .Z(clknet_leaf_94_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_95_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_95_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_96_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_96_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_97_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_97_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_98_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_98_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_99_wb_clk_i (.I(clknet_4_10__leaf_wb_clk_i),
    .Z(clknet_leaf_99_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_9_wb_clk_i (.I(clknet_4_4__leaf_wb_clk_i),
    .Z(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout100 (.I(net30),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 fanout101 (.I(net53),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout86 (.I(net87),
    .Z(net86));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout87 (.I(net88),
    .Z(net87));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout88 (.I(net89),
    .Z(net88));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout89 (.I(net15),
    .Z(net89));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 fanout90 (.I(net48),
    .Z(net90));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 fanout91 (.I(net67),
    .Z(net91));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 fanout92 (.I(net65),
    .Z(net92));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 fanout93 (.I(net63),
    .Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout94 (.I(net27),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout95 (.I(net42),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout96 (.I(net40),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout97 (.I(net34),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 fanout98 (.I(net33),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 fanout99 (.I(net32),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input1 (.I(io_in[10]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input10 (.I(io_in[7]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input11 (.I(io_in[8]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__buf_4 input12 (.I(io_in[9]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input2 (.I(io_in[11]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input3 (.I(io_in[12]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input4 (.I(io_in[13]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input5 (.I(io_in[33]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input6 (.I(io_in[34]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 input7 (.I(io_in[35]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 input8 (.I(io_in[5]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input9 (.I(io_in[6]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 max_cap85 (.I(_02766_),
    .Z(net85));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output13 (.I(net13),
    .Z(io_oeb[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output14 (.I(net14),
    .Z(io_oeb[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output15 (.I(net88),
    .Z(io_oeb[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output16 (.I(net16),
    .Z(io_oeb[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output17 (.I(net17),
    .Z(io_oeb[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output18 (.I(net18),
    .Z(io_oeb[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output19 (.I(net19),
    .Z(io_oeb[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output20 (.I(net20),
    .Z(io_oeb[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output21 (.I(net21),
    .Z(io_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output22 (.I(net22),
    .Z(io_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output23 (.I(net23),
    .Z(io_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output24 (.I(net24),
    .Z(io_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output25 (.I(net25),
    .Z(io_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output26 (.I(net26),
    .Z(io_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output27 (.I(net27),
    .Z(io_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output28 (.I(net28),
    .Z(io_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output29 (.I(net29),
    .Z(io_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output30 (.I(net30),
    .Z(io_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output31 (.I(net31),
    .Z(io_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output32 (.I(net32),
    .Z(io_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output33 (.I(net33),
    .Z(io_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output34 (.I(net34),
    .Z(io_out[24]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output35 (.I(net35),
    .Z(io_out[25]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output36 (.I(net36),
    .Z(io_out[26]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output37 (.I(net37),
    .Z(io_out[27]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output38 (.I(net38),
    .Z(io_out[28]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output39 (.I(net39),
    .Z(io_out[29]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output40 (.I(net40),
    .Z(io_out[30]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output41 (.I(net41),
    .Z(io_out[31]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output42 (.I(net42),
    .Z(io_out[32]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output43 (.I(net43),
    .Z(io_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output44 (.I(net44),
    .Z(io_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output45 (.I(net45),
    .Z(io_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output46 (.I(net46),
    .Z(io_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output47 (.I(net47),
    .Z(io_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output48 (.I(net90),
    .Z(la_data_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output49 (.I(net49),
    .Z(la_data_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output50 (.I(net50),
    .Z(la_data_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output51 (.I(net51),
    .Z(la_data_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output52 (.I(net52),
    .Z(la_data_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output53 (.I(net101),
    .Z(la_data_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output54 (.I(net54),
    .Z(la_data_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output55 (.I(net55),
    .Z(la_data_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output56 (.I(net56),
    .Z(la_data_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output57 (.I(net57),
    .Z(la_data_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output58 (.I(net58),
    .Z(la_data_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output59 (.I(net59),
    .Z(la_data_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output60 (.I(net60),
    .Z(la_data_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output61 (.I(net61),
    .Z(la_data_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output62 (.I(net62),
    .Z(la_data_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output63 (.I(net93),
    .Z(la_data_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output64 (.I(net64),
    .Z(la_data_out[24]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output65 (.I(net92),
    .Z(la_data_out[25]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output66 (.I(net66),
    .Z(la_data_out[26]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output67 (.I(net91),
    .Z(la_data_out[27]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output68 (.I(net68),
    .Z(la_data_out[28]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output69 (.I(net69),
    .Z(la_data_out[29]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output70 (.I(net70),
    .Z(la_data_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output71 (.I(net71),
    .Z(la_data_out[30]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output72 (.I(net72),
    .Z(la_data_out[31]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output73 (.I(net73),
    .Z(la_data_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output74 (.I(net74),
    .Z(la_data_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output75 (.I(net75),
    .Z(la_data_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output76 (.I(net76),
    .Z(la_data_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output77 (.I(net77),
    .Z(la_data_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output78 (.I(net78),
    .Z(la_data_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output79 (.I(net79),
    .Z(la_data_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 wire80 (.I(_01304_),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 wire81 (.I(_01188_),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 wire82 (.I(_01139_),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 wire83 (.I(_03694_),
    .Z(net83));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 wire84 (.I(_05750_),
    .Z(net84));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_102 (.ZN(net102));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_103 (.ZN(net103));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_104 (.ZN(net104));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_105 (.ZN(net105));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_106 (.ZN(net106));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_107 (.ZN(net107));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_108 (.ZN(net108));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_109 (.ZN(net109));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_110 (.ZN(net110));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_111 (.ZN(net111));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_112 (.ZN(net112));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_113 (.ZN(net113));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_114 (.ZN(net114));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_115 (.ZN(net115));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_116 (.ZN(net116));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_117 (.ZN(net117));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_118 (.ZN(net118));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_119 (.ZN(net119));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_120 (.ZN(net120));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_121 (.ZN(net121));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_122 (.ZN(net122));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_123 (.ZN(net123));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_124 (.ZN(net124));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_125 (.ZN(net125));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_126 (.ZN(net126));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_127 (.ZN(net127));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_128 (.ZN(net128));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_129 (.ZN(net129));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_130 (.ZN(net130));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_131 (.ZN(net131));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_132 (.ZN(net132));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_133 (.ZN(net133));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_134 (.ZN(net134));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_135 (.ZN(net135));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_136 (.ZN(net136));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_137 (.ZN(net137));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_138 (.ZN(net138));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_139 (.ZN(net139));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_140 (.ZN(net140));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_141 (.ZN(net141));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_142 (.ZN(net142));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_143 (.ZN(net143));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_144 (.ZN(net144));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_145 (.ZN(net145));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_146 (.ZN(net146));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_147 (.ZN(net147));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_148 (.Z(net148));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_149 (.Z(net149));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_150 (.Z(net150));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_151 (.Z(net151));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_152 (.Z(net152));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_153 (.Z(net153));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_154 (.Z(net154));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_155 (.Z(net155));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_156 (.Z(net156));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_157 (.Z(net157));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_158 (.Z(net158));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_159 (.Z(net159));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_160 (.Z(net160));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_161 (.Z(net161));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_162 (.Z(net162));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_163 (.Z(net163));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_164 (.Z(net164));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_165 (.Z(net165));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_166 (.Z(net166));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_167 (.Z(net167));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_168 (.Z(net168));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_169 (.Z(net169));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_170 (.Z(net170));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_171 (.Z(net171));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_172 (.Z(net172));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_173 (.Z(net173));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_174 (.Z(net174));
 assign io_oeb[0] = net148;
 assign io_oeb[13] = net153;
 assign io_oeb[14] = net102;
 assign io_oeb[15] = net103;
 assign io_oeb[16] = net104;
 assign io_oeb[17] = net105;
 assign io_oeb[18] = net106;
 assign io_oeb[19] = net107;
 assign io_oeb[1] = net149;
 assign io_oeb[20] = net108;
 assign io_oeb[21] = net109;
 assign io_oeb[22] = net110;
 assign io_oeb[23] = net111;
 assign io_oeb[24] = net112;
 assign io_oeb[25] = net113;
 assign io_oeb[26] = net114;
 assign io_oeb[27] = net115;
 assign io_oeb[28] = net116;
 assign io_oeb[29] = net117;
 assign io_oeb[2] = net150;
 assign io_oeb[30] = net118;
 assign io_oeb[31] = net119;
 assign io_oeb[32] = net120;
 assign io_oeb[33] = net154;
 assign io_oeb[34] = net155;
 assign io_oeb[35] = net156;
 assign io_oeb[36] = net157;
 assign io_oeb[37] = net158;
 assign io_oeb[3] = net151;
 assign io_oeb[4] = net152;
 assign io_out[0] = net121;
 assign io_out[13] = net126;
 assign io_out[1] = net122;
 assign io_out[2] = net123;
 assign io_out[33] = net127;
 assign io_out[34] = net128;
 assign io_out[35] = net129;
 assign io_out[36] = net130;
 assign io_out[37] = net131;
 assign io_out[3] = net124;
 assign io_out[4] = net125;
 assign la_data_out[32] = net159;
 assign la_data_out[33] = net132;
 assign la_data_out[34] = net160;
 assign la_data_out[35] = net133;
 assign la_data_out[36] = net161;
 assign la_data_out[37] = net134;
 assign la_data_out[38] = net162;
 assign la_data_out[39] = net135;
 assign la_data_out[40] = net163;
 assign la_data_out[41] = net136;
 assign la_data_out[42] = net164;
 assign la_data_out[43] = net137;
 assign la_data_out[44] = net165;
 assign la_data_out[45] = net138;
 assign la_data_out[46] = net166;
 assign la_data_out[47] = net139;
 assign la_data_out[48] = net140;
 assign la_data_out[49] = net167;
 assign la_data_out[50] = net141;
 assign la_data_out[51] = net168;
 assign la_data_out[52] = net142;
 assign la_data_out[53] = net169;
 assign la_data_out[54] = net143;
 assign la_data_out[55] = net170;
 assign la_data_out[56] = net144;
 assign la_data_out[57] = net171;
 assign la_data_out[58] = net145;
 assign la_data_out[59] = net172;
 assign la_data_out[60] = net146;
 assign la_data_out[61] = net173;
 assign la_data_out[62] = net147;
 assign la_data_out[63] = net174;
endmodule

