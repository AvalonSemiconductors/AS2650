* NGSPICE file created from wrapped_as2650.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_2 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_4 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyd_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyd_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai33_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai33_1 A1 A2 A3 B1 B2 B3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

.subckt wrapped_as2650 io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ vdd vss wb_clk_i
XFILLER_95_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7406__A1 _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6209__A2 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7963_ _1517_ _3088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_54_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6425__I _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6914_ _2105_ _2120_ _2121_ _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7894_ as2650.addr_buff\[0\] as2650.addr_buff\[1\] as2650.addr_buff\[2\] _3021_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_39_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4640__A1 _4212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6845_ _2030_ _2043_ _2056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8382__A2 _2215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6776_ _1958_ _1974_ _1988_ _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6393__A1 _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8515_ _2899_ _3610_ _3611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_52_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5727_ as2650.stack\[6\]\[14\] _0962_ _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_109_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4943__A2 _4140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8446_ _3164_ _3536_ _3543_ _3544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5658_ _0953_ _0903_ _0954_ _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6696__A2 _1909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4609_ as2650.ins_reg\[2\] as2650.ins_reg\[3\] _4190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_8377_ _2482_ _2354_ _3473_ _3476_ _3477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_102_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5589_ _4251_ _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_11_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7328_ _1308_ _2467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7205__B _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8087__I _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7259_ _1319_ _1347_ _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_46_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7948__A2 _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output37_I net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6620__A2 _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4631__A1 _4206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8373__A2 _3464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4934__A2 _4306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6136__A1 _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7884__A1 _2521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4698__A1 _4277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7636__A1 _2197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6439__A2 _4431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5414__I _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5111__A2 _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7769__C _2502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_60_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_60_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_67_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7939__A2 _3056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8061__A1 _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4960_ _4364_ _4514_ _4539_ _4363_ _4540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_52_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4891_ _4455_ _4462_ _4471_ _4472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_36_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8364__A2 _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6630_ _1795_ _1859_ _1860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_60_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6375__A1 _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6561_ as2650.r123_2\[1\]\[4\] _1719_ _1741_ _1792_ _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8116__A2 _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8300_ _2581_ _4380_ _3402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_121_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5512_ _0804_ _0808_ _0812_ _0816_ _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_9280_ _0173_ clknet_leaf_26_wb_clk_i net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__9305__CLK clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6492_ as2650.r123_2\[1\]\[0\] _1719_ _1724_ _1727_ _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_121_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8231_ _0910_ _2144_ _3334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7875__A1 _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5443_ _0748_ _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6678__A2 _1905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4689__A1 _4247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8162_ _1711_ _3266_ _3267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5350__A2 _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5374_ _0680_ _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7113_ _2278_ _2279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8093_ _3186_ _3204_ _1576_ _3205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7044_ _2233_ _2234_ _0121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_41_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7679__C _2565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8052__A1 _2535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8995_ _1287_ _4033_ _4034_ _0526_ _3199_ _4035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_103_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7946_ _4237_ _2348_ _3070_ _3071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_103_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7877_ _2991_ _3004_ _3005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5994__I _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8355__A2 _3423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6828_ _2035_ _2038_ _2039_ _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__5169__A2 _4386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4916__A2 _4414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6759_ _1964_ _1968_ _1972_ _1973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_17_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8658__A3 _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7866__A1 _2719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8429_ _3379_ _3495_ _3517_ _3527_ _3373_ _3528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_136_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5341__A2 _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7618__A1 _2719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5234__I _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4852__A1 _4427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8043__A1 _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4604__A1 _4181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5652__I0 _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8346__A2 _1919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9328__CLK clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5409__I as2650.r123\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6949__B _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7321__A3 _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7609__A1 _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5090_ _0354_ _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_42_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4983__I _4248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4843__A1 _4312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7800_ _2919_ _2505_ _2688_ _2362_ _2930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_80_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8780_ _1226_ _3793_ _3863_ _3864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_92_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5399__A2 _4481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5992_ _1260_ _1265_ _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_91_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7731_ _2824_ _2862_ _2863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4943_ _4520_ _4140_ _4521_ _4522_ _4523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_36_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6703__I _1923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7662_ _2782_ _2792_ _2794_ _2795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4874_ as2650.stack\[3\]\[8\] _4452_ _4454_ _4455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6613_ _4382_ _4284_ _1810_ _1841_ _1843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_18_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7593_ _2726_ _2727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6544_ _1757_ _1763_ _1776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9332_ _0225_ clknet_leaf_80_wb_clk_i as2650.r0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5571__A2 _4193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7848__A1 _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9263_ _0156_ clknet_leaf_52_wb_clk_i as2650.stack\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6475_ _4328_ _1688_ _1704_ _1711_ _1712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_12_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8214_ as2650.stack\[7\]\[0\] _1919_ _1638_ as2650.stack\[6\]\[0\] _3318_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_133_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5426_ _4427_ _0679_ _0731_ _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_133_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9194_ _0087_ clknet_leaf_48_wb_clk_i as2650.stack\[1\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6520__B2 _1753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8145_ as2650.cycle\[5\] _3243_ as2650.cycle\[3\] _3232_ _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_86_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5357_ _0349_ _4505_ _0369_ _0541_ _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_88_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5054__I _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8273__A1 _3055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7076__A2 _2256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8076_ _1391_ _3189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_141_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5288_ _0595_ _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7027_ _2223_ _4482_ _0968_ _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_59_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8576__A2 _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6587__A1 _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8978_ _4017_ _1467_ _4018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5938__B _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7929_ _2422_ _2453_ _3055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__8328__A2 _3355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6339__A1 _4316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5011__A1 _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7444__I net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7303__A3 _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7067__A2 _2248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5078__A1 _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8016__A1 _3120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8567__A2 _3481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9150__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7619__I _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5002__A1 _4277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8878__C _3923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4590_ _4162_ _4170_ _4171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9055__B _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6260_ _1517_ _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6502__A1 _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5305__A2 _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6502__B2 _4441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5211_ _4269_ _0519_ _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6191_ _0600_ _0821_ _1428_ _1448_ _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_48_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5142_ _0413_ _4331_ _0450_ _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5069__A1 _4399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8185__I _3288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6805__A2 _2017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5073_ _0361_ _4363_ _4408_ _0382_ _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_111_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8007__A1 _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8901_ _3958_ _3959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_49_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6281__A3 _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8558__A2 _3644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8832_ _2223_ _0624_ _0968_ _3912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_20_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6033__A3 _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8763_ _3844_ _2027_ _3846_ _3847_ _3810_ _3848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5975_ _1248_ _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7714_ _2837_ _2841_ _2845_ _2818_ _2846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_100_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4926_ _4505_ _4506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4595__A3 _4175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5792__A2 _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8694_ _3762_ _3763_ _3764_ _3782_ _3783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_139_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7645_ net34 _2778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4857_ _4202_ _4438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5049__I _4520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7576_ _2663_ _2710_ _2711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6741__A1 _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4788_ _4298_ _4369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9315_ _0208_ clknet_leaf_24_wb_clk_i as2650.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6527_ _1759_ _1731_ _1760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8494__A1 _3333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7297__A2 _2435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9246_ _0139_ clknet_leaf_62_wb_clk_i as2650.r123\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6458_ _1697_ _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5409_ as2650.r123\[0\]\[6\] _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_9177_ _0070_ clknet_leaf_71_wb_clk_i as2650.ins_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6389_ as2650.stack\[3\]\[8\] _1644_ _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_138_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8128_ _3179_ _3233_ _3238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8246__A1 _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8309__B _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8797__A2 _3557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8059_ _3168_ _3171_ _3172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9173__CLK clknet_leaf_60_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8549__A2 _3621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8823__I _3903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7439__I _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5783__A2 _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8979__B _1716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7883__B _2943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8021__I1 _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8721__A2 _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5535__A2 _4334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8485__A1 _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7288__A2 _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5838__A3 _4444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8237__A1 _4530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5471__A1 as2650.stack\[4\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5471__B2 as2650.stack\[5\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5223__B2 as2650.stack\[6\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5760_ _4210_ _1040_ _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4711_ _4291_ _4190_ _4292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5691_ _0961_ _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7430_ _0862_ _4390_ _2568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8712__A2 _4535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4642_ _4162_ _4223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_129_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5526__A2 _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6723__A1 _1934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7361_ _2499_ _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4573_ _4143_ _4153_ _4154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_128_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6312_ _1462_ _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9100_ _4122_ _4129_ _4130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8476__A1 _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7292_ _1163_ _2408_ _2406_ _2431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_9031_ _2450_ _3074_ _4067_ _4068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6243_ _0884_ _4167_ _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__7812__I _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9196__CLK clknet_leaf_47_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8228__A1 _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6174_ _4303_ _0403_ _0404_ _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_44_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8779__A2 _3792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6428__I _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5125_ _4477_ _0433_ _0434_ _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5332__I _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5056_ as2650.r123\[2\]\[3\] as2650.r123_2\[2\]\[3\] _4516_ _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_73_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5462__A1 _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8400__A1 _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6006__A3 _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8815_ _0834_ _2753_ _3889_ _3896_ _3897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_26_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8746_ _3810_ _0400_ _3831_ _1535_ _3832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_41_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5765__A2 _4261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5958_ _1230_ _1231_ _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8799__B _3780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4909_ _4487_ _4489_ _4490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5889_ _0592_ _1068_ _1069_ _1166_ _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_8677_ _3765_ _3766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8703__A2 _3368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7628_ _2727_ _2761_ _2762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_142_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6714__A1 as2650.stack\[0\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7559_ _0594_ _2694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6190__A2 _1447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8467__A1 _2825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9229_ _0122_ clknet_leaf_62_wb_clk_i as2650.r123_2\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7722__I _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8219__A1 as2650.stack\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6338__I as2650.psl\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5242__I _4332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5205__A1 _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6073__I _4167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6953__A1 _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5756__A2 _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4803__I1 as2650.r123\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7902__B1 _3028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_14_wb_clk_i clknet_3_2_0_wb_clk_i clknet_leaf_14_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_61_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6181__A2 _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8458__A1 _4477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6469__B1 _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5152__I as2650.holding_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7433__A2 _2569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8630__A1 _3329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6930_ _1223_ _1940_ _2019_ as2650.r123_2\[2\]\[7\] _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_81_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7197__A1 _4393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6861_ _2028_ _2071_ _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_62_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8600_ _2353_ _3691_ _3692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8933__A2 _3964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5812_ as2650.r123_2\[0\]\[1\] _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6792_ _1965_ _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8531_ _2333_ _3610_ _3626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5743_ _1000_ _1022_ _1028_ _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_37_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8462_ _2201_ _3377_ _1566_ _3560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5674_ _4487_ _0854_ _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7413_ _1569_ _2551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_11_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4707__B1 _4286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4625_ _4199_ _4205_ _4206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_8393_ _3492_ _3457_ _3288_ _3493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6172__A2 _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8449__A1 _3458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7344_ _1463_ _2482_ _2483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8449__B2 _3126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4556_ _4136_ _4137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4722__A3 _4302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5771__B _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7275_ _4209_ _2413_ _2414_ _1566_ _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_1_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9014_ _0621_ _4030_ _3216_ _4052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6226_ _1479_ _4187_ _1480_ _1481_ _1483_ _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XANTENNA__7672__A2 _2553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5683__A1 _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6157_ as2650.stack\[4\]\[9\] _1420_ _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5062__I _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5108_ _4330_ _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8621__A1 _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7424__A2 _4513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6227__A3 _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6088_ _1360_ _1227_ _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5997__I _4543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5435__A1 _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5039_ _4518_ _4523_ _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9211__CLK clknet_leaf_76_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8385__B1 _3322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8924__A2 _1823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8385__C2 as2650.stack\[5\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5738__A2 _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6935__A1 _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8729_ _3810_ _4388_ _3811_ _3815_ _3816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_142_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9361__CLK clknet_leaf_74_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8152__A3 _2719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7360__A1 _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7880__C _2852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput20 net20 io_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_134_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput31 net31 io_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput42 net42 io_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__5123__B1 _4470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6068__I _4263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6218__A3 _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5426__A1 _4427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7179__A1 _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8915__A2 _1753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6926__A1 _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5729__A2 _4466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6531__I _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7351__A1 _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8694__A4 _3782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5390_ _0571_ _0665_ _0663_ _4358_ _0487_ _0591_ _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__5901__A2 _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4986__I as2650.holding_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7060_ _2242_ _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7654__A2 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6457__A3 _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6011_ _1270_ _1274_ _1284_ _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_86_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7406__A2 _4528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8603__A1 _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6209__A3 _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8603__B2 _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9234__CLK clknet_leaf_62_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5610__I _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7962_ _2463_ _3086_ _3087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6090__A1 _4550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6913_ _2103_ _2116_ _2121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7030__C _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7893_ as2650.addr_buff\[4\] _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_23_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4640__A2 _4220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6844_ _2033_ _2054_ _2055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9384__CLK clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7590__A1 _2687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8119__B1 _3225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6775_ _1960_ _1973_ _1988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6393__A2 _1643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8514_ _0896_ _3609_ _3610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5726_ _1015_ _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8445_ _1526_ _2777_ _3541_ _3542_ _3070_ _3543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_5657_ as2650.stack\[5\]\[7\] _0904_ _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8796__C _3777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4608_ _4161_ _4171_ _4188_ _4189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8376_ _3082_ _3456_ _3475_ _3476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5588_ _0836_ _0880_ _0890_ _0891_ _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_89_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4896__I _4476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7327_ _2465_ _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8842__A1 _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7258_ _1571_ _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6209_ _1465_ _1232_ _1466_ _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_131_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7189_ _2335_ _2338_ _1324_ _1313_ _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7948__A3 _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4631__A2 _4211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7030__B1 _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8052__B _3164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7581__A1 _2181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5395__C _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8987__B _4026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6136__A2 _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5895__A1 _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4698__A2 _4278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9086__A1 _4041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7636__A2 _2580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8833__A1 _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9257__CLK clknet_leaf_55_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4870__A2 _4450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6526__I as2650.r0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8061__A2 _3153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8349__B1 _1638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8741__I _4365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9010__A1 _3214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4890_ as2650.stack\[0\]\[8\] _4466_ _4470_ as2650.stack\[1\]\[8\] _4471_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_83_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5586__B _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7572__A1 _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6375__A2 _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7572__B2 _2672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6261__I _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6560_ _1791_ _1792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_125_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5511_ _0651_ _0815_ _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6491_ _1726_ _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6127__A2 _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8667__A4 _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8230_ _3291_ _3333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5442_ _0610_ _0678_ _0743_ _0611_ _0747_ _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__6678__A3 _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4689__A2 _4262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5886__A1 _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8188__I _3291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5373_ _0679_ _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8161_ _3265_ _1527_ _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5605__I _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7112_ _2277_ _2278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7627__A2 _2697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8092_ _3136_ _3061_ _3176_ _3203_ _3204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_113_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8824__A1 _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8285__C1 as2650.stack\[5\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7025__C _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7043_ _0951_ _2224_ _2234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_87_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8137__B _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8588__B1 _3317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6436__I _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8052__A2 _3162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8994_ _1087_ _1287_ _4034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7976__B _2403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7945_ _2347_ _3070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4613__A2 _4192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9001__A1 _4479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7876_ _2960_ _2975_ _3004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6827_ _0585_ _1810_ _2039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7267__I _2406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5169__A3 _4524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6610__I0 as2650.r123\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6171__I _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6758_ _1966_ _1969_ _1971_ _1972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_109_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5709_ _0963_ _1000_ _1001_ _0019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7315__A1 _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6689_ as2650.stack\[1\]\[11\] _1911_ _1914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_87_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8428_ _3336_ _3496_ _3525_ _3369_ _3526_ _3527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__7866__A2 _2993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5877__A1 _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9068__A1 _3812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8359_ _3394_ _3459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8815__A1 _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5629__A1 _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8579__B1 _3670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4852__A2 _4430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8043__A2 _3155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4604__A2 _4184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5014__C1 _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6109__A2 _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7306__A1 _2436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8510__B _3604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7857__A2 _2950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9059__A1 _4316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7609__A2 _2703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8806__A1 _2635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8282__A2 _3322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5096__A2 _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4843__A2 _4423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8034__A2 _3148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5160__I _4191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6045__A1 _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5991_ _1261_ _1264_ _1233_ _1228_ _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_75_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7730_ _2751_ _2846_ _2861_ _2862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_79_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4942_ as2650.r123\[1\]\[2\] as2650.r123\[0\]\[2\] as2650.r123_2\[1\]\[2\] as2650.r123_2\[0\]\[2\]
+ _4139_ _4379_ _4522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__8404__C _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7661_ _2793_ _2794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4873_ _4453_ _4454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6612_ as2650.r0\[0\] _1841_ _1842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7592_ _0939_ net1 _2726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_127_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5020__A2 _4452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9331_ _0224_ clknet_leaf_80_wb_clk_i as2650.r0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6543_ _1768_ _1767_ _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_105_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7848__A2 _2976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9262_ _0155_ clknet_leaf_51_wb_clk_i as2650.stack\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6474_ _1710_ _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5859__A1 _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8213_ _2387_ _3317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5425_ _0730_ _0469_ _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9193_ _0086_ clknet_leaf_48_wb_clk_i as2650.stack\[1\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6520__A2 _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8144_ _2150_ _3250_ _1339_ _3178_ _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5356_ _0589_ _0574_ _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_134_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5287_ _0594_ _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8075_ _1570_ _3174_ _3185_ _3187_ _2400_ _3188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_101_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6284__A1 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7026_ _0957_ _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6284__B2 _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8576__A3 _3021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8977_ _1250_ _3773_ _4017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6587__A2 _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8981__B1 _2408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8381__I _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7928_ _1353_ _3050_ _3052_ _3053_ _3054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA__8314__C _2856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7859_ _2369_ _2985_ _2986_ _2987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7536__A1 _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6339__A2 _4391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5011__A2 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4770__A1 _4348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5245__I _4336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8264__A2 _3366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_39_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_39_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_120_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5078__A2 _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6275__A1 _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8016__A2 _3133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7775__A1 _2901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8291__I _3392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4589__A1 _4167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7527__A1 _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5002__A2 _4329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4761__A1 _4341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8488__C1 as2650.stack\[5\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6502__A2 _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5210_ _0492_ _4545_ _0515_ _0518_ _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_48_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6190_ _1444_ _1447_ _1448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8466__I _3562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5141_ _4257_ _4525_ _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8255__A2 _3335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7370__I _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5069__A2 _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5072_ _4538_ _4388_ _0381_ _4362_ _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_84_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8900_ _1601_ _4272_ _3958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8007__A2 _3126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8831_ _2285_ _3908_ _3909_ as2650.stack\[6\]\[1\] _3910_ _3911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_65_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8415__B _3510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6033__A4 _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8762_ _4434_ _3847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5974_ _1247_ _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7713_ _2842_ _2844_ _2845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_40_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4925_ _4283_ _4289_ _4381_ _4385_ _4505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_8693_ _1691_ _3766_ _2629_ _3781_ _3782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7518__B2 _2502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7644_ _2776_ _2777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4856_ _4436_ _4437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8191__A1 _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7575_ _2584_ _2585_ _2666_ _2664_ _2710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__7545__I _2403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4787_ _4367_ _4142_ _4368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6741__A2 _1732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9314_ _0207_ clknet_leaf_9_wb_clk_i as2650.psu\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6526_ as2650.r0\[2\] _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9245_ _0138_ clknet_3_0_0_wb_clk_i as2650.r123\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6457_ _1678_ _1354_ _0852_ _1346_ _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA__5065__I _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5408_ _0635_ _4440_ _0714_ _0005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_9176_ _0069_ clknet_leaf_59_wb_clk_i as2650.stack\[2\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6388_ _1642_ _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8127_ _3081_ _3236_ _3237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8246__A2 _2545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5339_ _0544_ _0645_ _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6257__A1 _1475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9318__CLK clknet_leaf_30_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8058_ _1249_ _3159_ _3169_ _3170_ _3171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_85_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7009_ _2206_ _2207_ _0113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8979__C _4018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4991__A1 as2650.holding_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8182__A1 _3052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8060__B _3172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4743__A1 _4323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8485__A2 _3574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5299__A2 _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8237__A2 _4380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7190__I _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5703__I _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6248__A1 _1492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7996__A1 _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5471__A2 _4481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7748__A1 _2866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8235__B _2926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8945__B1 _3993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5223__A2 _4478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6420__A1 as2650.stack\[2\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4710_ as2650.holding_reg\[0\] _4291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5690_ _0984_ _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8173__A1 _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4641_ _4221_ _4222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7920__A1 _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4734__A1 _4312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7360_ _0872_ _2151_ _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4572_ _4150_ _4152_ _4153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6202__C _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6311_ _4258_ _1212_ _1444_ _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8476__A2 _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7291_ _1939_ _2429_ _1347_ _2430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_144_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9030_ _3827_ _0516_ _2631_ _1034_ _4067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6242_ _4208_ _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8228__A2 _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6173_ _0813_ _1429_ _1430_ _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_135_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5124_ as2650.stack\[7\]\[10\] _0326_ _0427_ as2650.stack\[6\]\[10\] _0434_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7033__C _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7987__A1 _4264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5055_ _0364_ _4141_ _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5462__A2 _4547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7739__A1 _2866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8814_ _2630_ _1548_ _3895_ _3896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8400__A2 _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5214__A2 _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8745_ _3826_ _3830_ _3777_ _3831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5957_ _4219_ _4227_ _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_94_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4973__A1 _4154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4908_ _4143_ _4488_ _4432_ _4489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_8676_ _4394_ _3765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5888_ _0596_ _1072_ _1162_ _1165_ _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__8164__A1 as2650.psu\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7627_ _2760_ _2697_ _2728_ _2761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4839_ _4143_ _4420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__7911__A1 _3035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7558_ _2687_ _2532_ _2502_ _2692_ _2693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_135_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6509_ _4541_ _1733_ _1743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8467__A2 _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7489_ _2615_ _2625_ _2573_ _2626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_49_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6478__A1 _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__9140__CLK clknet_leaf_46_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9228_ _0121_ clknet_leaf_40_wb_clk_i as2650.stack\[4\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5150__A1 _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5150__B2 _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9159_ _0052_ clknet_leaf_58_wb_clk_i as2650.stack\[4\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8219__A2 _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5523__I _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7978__A1 _3087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6354__I as2650.psl\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_6_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6402__A1 as2650.stack\[3\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5205__A2 _4399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4803__I2 as2650.r123_2\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4964__A1 _4422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8155__A1 _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7902__A1 _2836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7185__I _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7902__B2 _2720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_54_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_4_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6469__A1 _4160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6469__B2 _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6529__I _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5141__A1 _4257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5692__A2 _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7969__A1 _3093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8630__A2 _3706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8918__B1 _3964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6860_ _2057_ _2070_ _2071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_74_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8394__A1 _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7197__A2 _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5811_ _1032_ _1055_ _1092_ _0030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6791_ _4519_ _1965_ _2004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8530_ _2382_ _3058_ _3625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5742_ as2650.stack\[5\]\[11\] _1025_ _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4955__A1 _4387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8146__A1 _2484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8461_ _3333_ _3530_ _3549_ _3558_ _3288_ _3559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5673_ _4152_ _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5608__I _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7412_ _2549_ _2550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4707__A1 _4285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4624_ _4149_ _4204_ _4205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__9163__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8392_ _2388_ _3492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4707__B2 _4287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7343_ _2481_ _2482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4555_ _4135_ _4136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5771__C _4438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7274_ net23 _2413_ _2414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9013_ _4050_ _3113_ _3114_ _1296_ _4051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_103_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6225_ _1482_ _1369_ _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_48_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5683__A2 _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6156_ _1415_ _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5107_ _4315_ _0406_ _0412_ _0416_ _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_57_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7698__C _2554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8621__A2 _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6087_ _4215_ _0874_ _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6632__A1 _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5435__A2 _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5499__B _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5038_ _0287_ _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6989_ _2190_ _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8728_ _3769_ _1749_ _3814_ _4435_ _1623_ _3815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_107_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8659_ _2927_ _3747_ _0971_ _3748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_103_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5371__A1 _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8829__I _3905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7648__B1 _2534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput21 net21 io_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput32 net32 io_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_107_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput43 net43 io_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_122_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5253__I _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5674__A2 _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6623__A1 _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5426__A2 _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8376__A1 _3082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7908__I as2650.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6926__A2 _2109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9186__CLK clknet_leaf_73_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8679__A2 _3326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7351__A2 _2478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7643__I _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8300__A1 _2581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6259__I _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6457__A4 _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5665__A2 _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6010_ _1277_ _1281_ _1233_ _1283_ _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_98_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input3_I io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5417__A2 _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7961_ _3072_ _3073_ _3079_ _3085_ _3086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_36_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6090__A2 _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6912_ _2103_ _2116_ _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7892_ net52 _2377_ _2852_ _3019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_82_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8367__A1 _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6843_ _2042_ _2054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_63_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4928__A1 _4282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8119__A1 _3208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6774_ _1956_ _1957_ _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_56_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7590__A2 _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8513_ _3607_ _3566_ _3608_ _3609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5725_ as2650.pc\[14\] _0858_ _0972_ as2650.r123_2\[0\]\[6\] _1014_ _1015_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_50_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8444_ _3537_ _3540_ _3181_ _3542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5656_ _0952_ _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5353__A1 _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4607_ _4176_ _4187_ _4188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8375_ _1582_ _2533_ _1508_ _3474_ _3475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__7553__I _2507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5587_ _0877_ _0870_ _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7326_ _2464_ _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_137_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7257_ _2394_ _2397_ _2398_ _1410_ _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_117_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6208_ _1320_ _1247_ _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7188_ _2337_ _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6139_ _1397_ _1405_ _1406_ _1392_ _0044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5801__I _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6605__A1 _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8333__B _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7030__A1 _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7030__B2 as2650.stack\[4\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7581__A2 _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8530__A1 _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5895__A2 _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4942__I1 as2650.r123\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8833__A2 _3912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5912__S _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8508__B _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9330__D _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8597__A1 _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6072__A2 _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9010__A2 _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7638__I _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7021__A1 _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7572__A2 _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5510_ _0813_ _0799_ _0814_ _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6490_ _1725_ _1718_ _1726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8521__A1 _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5441_ _0348_ _0746_ _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4689__A3 _4269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5886__A2 _4420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8160_ _4420_ _3265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__9077__A2 _4110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5372_ _0678_ _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_86_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7111_ _0622_ _2208_ _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7088__A1 _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9201__CLK clknet_leaf_60_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8285__B1 _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8091_ _2888_ _3202_ _3203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8285__C2 _1654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8824__A2 _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7042_ _2205_ _2219_ _2220_ as2650.stack\[4\]\[7\] _2209_ _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_86_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8588__A1 _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8588__B2 _3665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9351__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8993_ _4010_ _4028_ _4032_ _4033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_94_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7260__A1 _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7944_ _2349_ _3068_ _3069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6653__S _4144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5810__A2 _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4613__A3 _4193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7875_ _1575_ _3002_ _3003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__9001__A2 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6826_ as2650.r0\[4\] _1841_ _2038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7563__A2 _2697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8760__A1 as2650.psu\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6610__I1 as2650.r123_2\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6757_ _4519_ _1970_ _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5708_ as2650.stack\[6\]\[11\] _0986_ _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6688_ _1666_ _1908_ _1913_ _0086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7315__A2 _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8427_ _3290_ _3526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5639_ _0937_ _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8358_ _3393_ _3458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__9068__A2 _4097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7079__A1 _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7079__B2 as2650.stack\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7309_ _1230_ _1471_ _1231_ _1368_ _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_65_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8289_ _3095_ _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8815__A2 _2753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6826__A1 as2650.r0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5629__A2 _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5185__S0 _4196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8328__B _2182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8579__A1 _3459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8579__B2 _3504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4852__A3 _4432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7251__A1 _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8063__B _2607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6362__I _1618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7003__A1 _2200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5014__B1 _4460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8751__A1 _3189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8503__A1 _2204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7306__A2 _2441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5317__A1 as2650.stack\[2\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8289__I _3095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9224__CLK clknet_leaf_39_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4610__I _4190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8267__B1 _3368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8806__A2 _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6817__A1 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9374__CLK clknet_leaf_77_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7490__A1 _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6045__A2 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8752__I _3763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5990_ _1263_ _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4941_ _4286_ _4521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7368__I _2506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6272__I _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7660_ _1271_ _2793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4872_ as2650.psu\[2\] _4449_ _4453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__8742__A1 as2650.psu\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6611_ _1840_ _1841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7591_ _2579_ _2724_ _2725_ _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_53_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8701__B _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9330_ _0223_ clknet_leaf_80_wb_clk_i as2650.r0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6542_ _1769_ _1767_ _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_9_wb_clk_i clknet_3_3_0_wb_clk_i clknet_leaf_9_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_9_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9261_ _0154_ clknet_leaf_54_wb_clk_i as2650.stack\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6473_ _1709_ _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5616__I _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8212_ _3214_ _3313_ _3315_ _3316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5859__A2 _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5424_ as2650.holding_reg\[6\] _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9192_ _0085_ clknet_leaf_48_wb_clk_i as2650.stack\[1\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_86_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8143_ _4171_ _3250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5355_ _0661_ _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8074_ _2421_ _3186_ _3187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5286_ net10 _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8273__A3 _3285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6284__A2 _1534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6447__I _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7025_ _2170_ _2219_ _2220_ as2650.stack\[4\]\[1\] _2221_ _2222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_60_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7233__A1 _4357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8976_ _1482_ _3163_ _0875_ _4016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_56_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7784__A2 _2895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8981__B2 _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5795__A1 _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7927_ _4491_ _2446_ _3053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7858_ _2880_ _2950_ _2744_ _2986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6115__C _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7536__A2 _2592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8733__A1 _3763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6809_ _1984_ _2016_ _2020_ _2021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_141_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9247__CLK clknet_leaf_62_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7789_ net37 _2919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4770__A2 _4350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8058__B _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6275__A2 _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6357__I _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7224__A1 _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8421__B1 _3362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8972__A1 _2926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7188__I _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7527__A2 _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5538__A1 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8521__B _3046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8488__B1 _3361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8488__C2 _3362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5140_ _0401_ _0399_ _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6267__I as2650.psl\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6510__I0 as2650.r123\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5071_ _4378_ _0372_ _0380_ _4222_ _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_42_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5474__B1 _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7215__A1 _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8830_ _3900_ _3910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8415__C _3513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8761_ _1033_ _3772_ _3845_ _3846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_64_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5973_ _0868_ _4423_ _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7712_ _2784_ _2816_ _2843_ _2844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4924_ _4305_ _4306_ _4503_ _4504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_8692_ _3767_ _1383_ _3779_ _3780_ _3781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_127_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8715__A1 _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7643_ _2503_ _2776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4855_ _4419_ _4435_ _4436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8191__A2 _2487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7574_ _1581_ _0578_ _2708_ _2709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_119_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4786_ _4366_ _4367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9313_ _0206_ clknet_leaf_18_wb_clk_i as2650.cycle\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6525_ _1757_ _1746_ _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9244_ _0137_ clknet_leaf_39_wb_clk_i as2650.stack\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6456_ _1695_ _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_109_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5407_ _4274_ _0703_ _0713_ _0538_ _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__5701__A1 _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9175_ _0068_ clknet_leaf_60_wb_clk_i as2650.stack\[2\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6387_ _1642_ _1643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8126_ _0869_ _2506_ _3236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5338_ _0642_ _0644_ _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_138_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7454__A1 _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8057_ _3045_ _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5269_ _0571_ _0572_ _0573_ _0576_ _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_60_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7008_ _0951_ _2176_ _2207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7206__A1 _2351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8392__I _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8403__B1 _3500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5768__A1 _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8959_ _4002_ _4003_ _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8706__A1 as2650.psl\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8341__B _3441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4991__A2 _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8182__A2 _3069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5940__A1 _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8995__C _3199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7445__A1 _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6248__A2 _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8642__B1 _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8642__C2 as2650.pc\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7996__A2 _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6815__I _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7748__A2 _2876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8945__A1 _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5759__A1 _4157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4982__A2 _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5367__S _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4640_ _4212_ _4220_ _4221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7920__A2 _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4571_ _4151_ _4152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5931__A1 _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4734__A2 _4314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6310_ _1564_ _1567_ _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7290_ _1095_ _1324_ _2429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6241_ _1498_ _1248_ _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6172_ _1429_ _0753_ _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5115__B _4454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5123_ as2650.stack\[4\]\[10\] _0429_ _4470_ as2650.stack\[5\]\[10\] _0433_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_112_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7987__A2 _2824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5054_ _0363_ _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6725__I _1716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7739__A2 _2867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8813_ _1577_ _3894_ _3895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8744_ _1235_ _1764_ _3829_ _4434_ _3830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_5956_ _4185_ _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_53_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4907_ _4191_ _4488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_94_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8675_ _4398_ _2632_ _3764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5887_ _1163_ _1164_ _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8164__A2 _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7626_ _0933_ _0594_ _2760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4838_ _4418_ _4419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7372__B1 _2508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7911__A2 _2495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7557_ _1582_ _2688_ _2691_ _2648_ _2692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_105_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4769_ _4349_ _4244_ _4350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6508_ _0359_ _1722_ _1742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7488_ _0921_ _2528_ _2623_ _2550_ _2624_ _2625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_119_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7675__A1 _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6478__A2 _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6439_ _1253_ _4431_ _1681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_9227_ _0120_ clknet_leaf_36_wb_clk_i as2650.stack\[4\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5804__I _4170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9158_ _0051_ clknet_leaf_56_wb_clk_i as2650.stack\[4\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5150__A2 _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5150__B3 _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8109_ _3219_ _3212_ _3220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9089_ _1319_ _2925_ _1245_ _4119_ _4120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_88_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_4_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5679__C _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4661__A1 _4235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4803__I3 as2650.r123_2\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4964__A2 _4194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5187__S _4516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8155__A2 _3257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6370__I _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6166__A1 _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7902__A2 _3026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9104__A1 _3133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7666__A1 _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6469__A2 _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5714__I _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9333__D _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4758__C _4338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7134__C _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5141__A2 _4525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7418__A1 _4390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7969__A2 _2155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_23_wb_clk_i clknet_3_3_0_wb_clk_i clknet_leaf_23_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8091__A1 _2888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8918__A1 _3962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8394__A2 _3374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5810_ _1056_ _1084_ _1091_ _1054_ _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6790_ _2000_ _2002_ _2003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_37_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5741_ _0993_ _1022_ _1027_ _0025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__9077__B _3619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4955__A2 _4534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8146__A2 _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8460_ _3216_ _3550_ _3557_ _3481_ _3371_ _3558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__9308__CLK clknet_leaf_18_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5672_ _0967_ _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7411_ _2523_ _2549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4623_ _4201_ _4203_ _4204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_8391_ _3210_ _3457_ _3490_ _3491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4707__A2 _4140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5904__A1 _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7342_ _0853_ _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4554_ as2650.ins_reg\[1\] _4135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5380__A2 _4193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7273_ _2403_ _2405_ _2412_ _2400_ _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__5624__I _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9012_ _0620_ _4030_ _4050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6224_ _0867_ _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7409__A1 _2530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6155_ _0976_ _1417_ _1419_ _0047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_112_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5106_ _0413_ _0414_ _4314_ _0415_ _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6086_ _1354_ _1356_ _1358_ _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8156__B _3229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6455__I _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6632__A2 _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5037_ as2650.r123\[0\]\[2\] _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5435__A3 _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7995__B _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8385__A2 _3319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6988_ _2189_ _2190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8603__C _2855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8727_ _3812_ _3772_ _3813_ _3814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5939_ _0834_ _1071_ _1213_ _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_55_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4703__I as2650.r0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6148__A1 net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8658_ _4160_ _3265_ _1288_ _3747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_142_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7896__A1 _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7609_ _0685_ _2703_ _2743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8589_ _3680_ _3681_ _3526_ _3682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_31_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7648__A1 _2778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7648__B2 _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput11 net11 io_oeb[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_108_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput22 net22 io_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput33 net33 io_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput44 net44 io_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_107_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5123__A2 _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6320__A1 _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7889__C _2961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8073__A1 _4417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7820__A1 _2662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6365__I _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6623__A2 _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8376__A2 _3456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9328__D _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7129__C _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5872__C _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8021__S _3130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7639__A1 _2757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5444__I _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8300__A2 _4380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6311__A1 _4258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8064__A1 _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7811__A1 _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7811__B2 _2940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7960_ _3080_ _3084_ _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4625__A1 _4199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6911_ _1201_ _1940_ _1942_ as2650.r123_2\[2\]\[6\] _2119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__9013__B1 _3114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7891_ _1711_ _3017_ _3018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8367__A2 _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6842_ _1994_ _2045_ _2053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_1_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9130__CLK clknet_leaf_58_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6773_ _1949_ _1976_ _1985_ _1986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4928__A2 _4288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8119__A2 _3209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8512_ _1616_ _4370_ _3608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5724_ _0715_ _4416_ _1009_ _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5655_ as2650.pc\[7\] _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8443_ _3537_ _3540_ _3541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__9280__CLK clknet_leaf_26_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4606_ as2650.ins_reg\[3\] _4186_ _4187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_8374_ as2650.addr_buff\[4\] _2754_ _3474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5586_ _0881_ _0882_ _0889_ _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6550__A1 _4285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7325_ _2426_ _2456_ _2463_ _2464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_11_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7256_ net24 _2394_ _2398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_46_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5105__A2 _4526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6302__A1 _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6207_ _1464_ _1355_ _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7187_ _2336_ _4241_ _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4864__A1 _4415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8055__A1 _3158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6138_ net19 _1402_ _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8055__B2 _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6185__I _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7802__A1 _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6069_ _1340_ _1341_ _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9004__B1 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6369__A1 _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8333__C _2651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7030__A2 _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5041__A1 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5529__I _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7869__A1 _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8530__A2 _3058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6541__A1 _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4855__A1 _4419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8046__A1 _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6309__B _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8597__A2 _3669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9153__CLK clknet_leaf_16_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4607__A1 _4176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8524__B _3619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8349__A2 _1919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7919__I _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7557__B1 _2691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9010__A3 _3126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5583__A2 _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6780__A1 _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8521__A2 _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5440_ _0745_ _0716_ _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_121_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6532__A1 _4405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5335__A2 _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5371_ _0673_ _0675_ _0677_ _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__5886__A3 _4204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7110_ _2276_ _0145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8090_ _3178_ _3192_ _3179_ _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_99_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8285__B2 as2650.stack\[4\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8824__A3 _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7041_ _2200_ _2211_ _2232_ _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_113_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8037__A1 _2416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8588__A2 _3327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8992_ _2794_ _0342_ _4031_ _4032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_94_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout54_I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7260__A2 _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7943_ _3065_ _3067_ _3068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7874_ _0997_ _2525_ _3000_ _3001_ _3002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_63_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_7_0_wb_clk_i clknet_0_wb_clk_i clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_6825_ _2034_ _2009_ _2036_ _2037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8760__A2 _3772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5574__A2 _4175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6756_ _1840_ _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6771__A1 _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5707_ _0999_ _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6687_ as2650.stack\[1\]\[10\] _1911_ _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8512__A2 _4370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7315__A3 _2351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8426_ _3521_ _3524_ _3525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5326__A2 _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5638_ _0711_ _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_30_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8357_ _3456_ _3457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5569_ _0867_ _0872_ _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5084__I _4278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7308_ _1087_ _2446_ _2447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8288_ _3383_ _3384_ _3385_ _3389_ _3390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_132_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7239_ _1252_ _2380_ _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5185__S1 _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5812__I as2650.r123_2\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9176__CLK clknet_leaf_59_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_69_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7251__A2 _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output35_I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8751__A2 _3836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5565__A2 _4369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8503__A2 _3570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7306__A3 _2442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5317__A2 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8267__A1 _3199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8267__B2 _3369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6817__A2 _2027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4828__A1 _4406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8019__A1 _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7490__A2 _2580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6981__C _2173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4940_ _4519_ _4520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_45_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4871_ _4451_ _4452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5005__A1 _4332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6610_ as2650.r123\[0\]\[6\] as2650.r123_2\[0\]\[6\] _4145_ _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7590_ _2687_ _2466_ _1635_ _2725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6541_ _1156_ _1715_ _1773_ _0079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7384__I _2517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6472_ _1708_ _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5308__A2 _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6505__A1 _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9260_ _0153_ clknet_leaf_50_wb_clk_i as2650.stack\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8211_ _2145_ _2794_ _3194_ _3314_ _3315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5423_ _0720_ _0727_ _0728_ _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_9191_ _0084_ clknet_leaf_47_wb_clk_i as2650.stack\[1\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9199__CLK clknet_leaf_47_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5354_ _0636_ _0641_ _0658_ _0660_ _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8142_ _1301_ _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8073_ _4417_ _1279_ _3186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5285_ _0592_ _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4819__A1 _4398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5632__I _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8148__C _3207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7024_ _2209_ _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5492__A1 _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7769__B1 _2535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8430__A1 _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7233__A2 _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8975_ _4014_ _4015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8164__B _3268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7559__I _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5244__A1 _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8981__A2 _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7926_ _2457_ _2425_ _3051_ _3052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_82_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7857_ _2953_ _2950_ _2612_ _2985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6808_ _1986_ _2015_ _2020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_7788_ _2476_ _2916_ _2917_ _2554_ _2918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8611__C _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6739_ as2650.r0\[5\] _1761_ _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5807__I _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8497__A1 _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8409_ _1180_ _0583_ _3507_ _3508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_9389_ _0282_ clknet_leaf_6_wb_clk_i as2650.psu\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8249__A1 _2335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8058__C _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8421__B2 as2650.stack\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8972__A2 _4011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8802__B _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_48_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8724__A2 _3390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5538__A2 _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9336__D _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4621__I net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8488__A1 as2650.stack\[7\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9341__CLK clknet_leaf_51_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7160__A1 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5452__I _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5070_ _0376_ _4397_ _0379_ _4230_ _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_69_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8660__A1 _4419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6510__I1 as2650.r123_2\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5474__A1 as2650.stack\[3\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7215__A2 _2363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8412__A1 _2196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8963__A2 _3989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8760_ as2650.psu\[4\] _3772_ _3845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5972_ _1229_ _1233_ _1245_ _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_80_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7711_ _0945_ net2 _2843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4923_ as2650.addr_buff\[6\] _4355_ _4503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_55_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8691_ _4394_ _3780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7642_ _0948_ _2655_ _2775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6726__A1 _1612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4854_ _4434_ _4435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7573_ _2706_ _2707_ _2708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4785_ as2650.r0\[7\] _4366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9312_ _0205_ clknet_leaf_18_wb_clk_i as2650.cycle\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8479__A1 _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6524_ as2650.r0\[1\] _1757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9243_ _0136_ clknet_leaf_55_wb_clk_i as2650.stack\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6455_ _0877_ _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5406_ _0438_ _0710_ _0712_ _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_9174_ _0067_ clknet_leaf_60_wb_clk_i as2650.stack\[2\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6386_ _1641_ _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5701__A2 _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8125_ _1451_ _3234_ _3235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5337_ _0543_ _0546_ _0643_ _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6458__I _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5362__I _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7454__A2 _2553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8651__A1 _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8056_ _1612_ _1256_ _1229_ _2482_ _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__6257__A3 _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5268_ _0384_ _0574_ _0575_ _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_9_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7007_ _2205_ _2171_ _2172_ as2650.stack\[2\]\[7\] _2141_ _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_60_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5199_ _0507_ _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8403__A1 _2996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6193__I _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9214__CLK clknet_leaf_41_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8958_ _3995_ _2117_ _4003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5768__A2 _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7909_ _2385_ _3028_ _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8889_ _1663_ _3948_ _3952_ _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_58_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8706__A2 _3792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6717__A1 _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9364__CLK clknet_leaf_73_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8341__C _2925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8182__A3 _3071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7390__A1 _2525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5940__A2 _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7142__A1 _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7142__B2 as2650.stack\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6350__C1 _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5272__I _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8642__A1 _4264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7445__A2 _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6248__A3 _1496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5456__A1 _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5208__A1 _4212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7748__A3 _2878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4616__I _4196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8945__A2 _3992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5759__A2 _4242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6708__A1 as2650.stack\[0\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7381__A1 _2416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5447__I _4376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4570_ as2650.halted net5 _4151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_50_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6240_ _1497_ _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7684__A2 _2816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8881__A1 _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6171_ _0548_ _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5182__I _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5122_ _0425_ _0428_ _0431_ _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7436__A2 _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8633__A1 _3703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6495__I0 as2650.r123\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9237__CLK clknet_leaf_55_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5053_ _0362_ _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7739__A3 _2869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8812_ _3890_ _3893_ _1629_ _3894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8743_ _3827_ _3773_ _3828_ _3829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5955_ _1228_ _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4906_ _4211_ _4487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8674_ _3757_ _3763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5886_ _1033_ _4420_ _4204_ _4211_ _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_107_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7625_ _2756_ _2749_ _2758_ _2759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4837_ _4417_ _4418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7372__A1 _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6175__A2 _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7372__B2 _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7556_ _2687_ _2690_ _2691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4768_ as2650.idx_ctrl\[1\] _4349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_5_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6507_ _1726_ _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7124__A1 _2285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7487_ _1569_ _2624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4699_ _4138_ as2650.ins_reg\[1\] _4280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_88_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9226_ _0119_ clknet_leaf_37_wb_clk_i as2650.stack\[4\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6438_ _1679_ _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7675__A2 _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8872__A1 _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8872__B2 as2650.stack\[7\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9157_ _0050_ clknet_leaf_57_wb_clk_i as2650.stack\[4\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6369_ _0790_ _1571_ _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8624__A1 _3093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8108_ _3158_ _3219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_62_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9088_ _1523_ _0339_ _4062_ _4119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_114_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5438__A1 _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8039_ _3151_ _1677_ _3152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5989__A2 _4330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4661__A2 _4241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8352__B _3420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5913__A2 _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9104__A2 _4028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7666__A2 _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8863__A1 _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7418__A2 _4352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5429__A1 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5429__B2 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8918__A2 _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_63_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_63_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__9040__A1 _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5601__A1 as2650.stack\[5\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5740_ as2650.stack\[5\]\[10\] _1025_ _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_37_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7354__A1 _2150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5177__I _4269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5671_ _0857_ _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7410_ _2529_ _2541_ _2547_ _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4622_ _4202_ _4203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8390_ _3480_ _3489_ _3490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5904__A2 _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4553_ net26 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7341_ _2479_ _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7272_ _2407_ _2408_ _1483_ _2409_ _2411_ _2412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_116_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9011_ _4026_ _4048_ _4049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6223_ _1320_ _1250_ _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_143_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7409__A2 _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8606__A1 _3046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6154_ as2650.stack\[4\]\[8\] _1418_ _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_140_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4891__A2 _4462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5105_ _0414_ _4526_ _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_131_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6085_ _4551_ _1357_ _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6093__A1 _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5036_ _4497_ _4499_ _0346_ _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_113_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9031__A1 _2450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7042__B1 _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6987_ _2188_ _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6471__I _1604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8726_ _0849_ _3773_ _3813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5938_ _0836_ _1072_ _1067_ _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8599__S _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8657_ _3743_ _3745_ _1516_ _3746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_139_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5869_ _1147_ _1146_ _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5087__I _4341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7608_ _1180_ _0698_ _2741_ _2742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_8588_ _0533_ _3327_ _3317_ _3665_ _3681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_124_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9098__A1 as2650.psu\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7539_ _2472_ _2674_ _2675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7648__A2 _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8845__A1 _2265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput12 net12 io_oeb[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput23 net23 io_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput34 net34 io_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_134_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9209_ _0102_ clknet_leaf_75_wb_clk_i as2650.r123_2\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4706__I0 as2650.r123\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput45 net45 io_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_89_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8073__A2 _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6084__A1 _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7820__A2 _2871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5831__A1 _4542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8861__I _3923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9022__A1 _2776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7033__B1 _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5595__B1 _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6139__A2 _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7336__A1 _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_117_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9089__A1 _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8836__A1 _2294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6311__A2 _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8257__B _4473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8064__A2 _3175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7272__B1 _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7811__A2 _2684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6910_ _1189_ _1937_ _2118_ _0103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9013__A1 _4050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8771__I _3757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7890_ _3012_ _3016_ _3017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_35_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6841_ _2026_ _2044_ _2052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7387__I _2524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7575__A1 _2584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6291__I _4391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6772_ _1952_ _1975_ _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4928__A3 _4381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8511_ _1616_ _4370_ _3607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5723_ _0977_ _1012_ _1013_ _0021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8720__B _3080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8442_ _3538_ _3507_ _3539_ _3540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_31_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5654_ _0791_ _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5889__A1 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4605_ _4179_ _4185_ _4186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8373_ _2353_ _3464_ _3473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5585_ _0883_ _0888_ _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6550__A2 _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8827__A1 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7324_ _2457_ _2462_ _2463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8946__I _3961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7255_ _1451_ _2396_ _1350_ _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_46_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6302__A2 _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6206_ _0884_ _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7186_ _1303_ _2336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_59_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8167__B _3151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4864__A2 _4444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6137_ _0711_ _1398_ _1404_ _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8055__A2 _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6066__A1 _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7802__A2 _2496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6068_ _4263_ _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5813__A1 _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5019_ as2650.stack\[7\]\[9\] _0326_ _0329_ _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__9004__A1 _4042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9004__B2 _3123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6369__A2 _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8763__B1 _3846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5041__A2 _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8709_ _1519_ _4514_ _1480_ _3797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_139_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7318__A1 _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7869__A2 _2984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6541__A2 _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8818__A1 _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4942__I3 as2650.r123_2\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8856__I _3928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8294__A2 _3355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8077__B _3189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4855__A2 _4435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8046__A2 _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6057__A1 _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5213__C _4262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4607__A2 _4187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7557__A1 _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7557__B2 _2648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9010__A4 _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7000__I _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8540__B _3095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7309__A1 _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7935__I _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6780__A2 _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6532__A2 _1764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8809__A1 _1611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5370_ _4300_ _0676_ _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5886__A4 _4211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8766__I _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8285__A2 _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5099__A2 _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7040_ _2201_ _2214_ _2217_ as2650.stack\[4\]\[6\] _2221_ _2232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__6286__I _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8037__A2 _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5190__I _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6048__A1 _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8991_ _4029_ _0360_ _4030_ _4031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7942_ _0891_ _3066_ _3067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7260__A3 _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7548__A1 _2579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7873_ _2149_ _3001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6235__B _4417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6824_ _1971_ _2035_ _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_1_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8006__I _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6220__A1 _4187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6755_ as2650.r0\[3\] _1810_ _1969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5706_ _0997_ _0980_ _0973_ as2650.r123_2\[0\]\[3\] _0998_ _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_108_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6686_ _1663_ _1908_ _1912_ _0085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_109_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8425_ _0525_ _3522_ _3523_ _3524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5637_ _0932_ _0861_ _0936_ _0012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7720__A1 _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5365__I _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8356_ _2188_ _3455_ _3456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5568_ _0868_ _0871_ _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7307_ _4422_ _4430_ _4432_ _1470_ _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__8676__I _4394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8287_ as2650.stack\[6\]\[2\] _3386_ _3388_ _3389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5499_ _0802_ _0803_ _0448_ _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_137_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7238_ _4179_ _1360_ _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_137_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7169_ _2294_ _2322_ _2325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6039__A1 _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7787__A1 _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8625__B _3500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7251__A3 _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8344__C _2856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7539__A1 _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5014__A2 _4481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6211__A1 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5565__A3 _4313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7306__A4 _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7711__A1 _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6278__A1 _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9120__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8019__A2 _3136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7778__A1 _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7778__B2 _2681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9270__CLK clknet_leaf_12_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4870_ _4448_ _4450_ _4451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5005__A2 _4386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6202__A1 _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7950__A1 _2450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6540_ as2650.r123_2\[1\]\[3\] _1719_ _1741_ _1772_ _1773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_53_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6471_ _1604_ _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7702__A1 _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6505__A2 _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8210_ _2335_ _3295_ _3314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5422_ _0719_ _0727_ _0411_ _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_9190_ _0083_ clknet_leaf_65_wb_clk_i as2650.r123_2\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5713__B1 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8141_ _2416_ _3248_ _0204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5353_ _0565_ _0659_ _0396_ _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_47_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8429__C _3373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4957__C _4231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8072_ _3177_ _3180_ _3184_ _3185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_88_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5284_ _0591_ _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4819__A2 _4399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7023_ _2216_ _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5492__A2 _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7769__A1 _2884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7769__B2 _2899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8430__A2 _3289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8974_ _3045_ _1246_ _1265_ _4013_ _3273_ _4014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_83_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6441__A1 _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5244__A2 _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7925_ _1480_ _2427_ _3051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7856_ _2982_ _2983_ _2984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_24_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8194__A1 _4392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6807_ _1941_ _2019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7787_ _2361_ _2870_ _2917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4999_ _4302_ _4326_ _0305_ _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_6738_ _1874_ _1950_ _1951_ _1886_ _1893_ _1952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_104_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8497__A2 _3374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6669_ _1865_ _1897_ _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8408_ _3505_ _3468_ _3506_ _3507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_30_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9143__CLK clknet_leaf_67_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9388_ _0281_ clknet_3_1_0_wb_clk_i net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8339_ _0508_ _0366_ _3439_ _3440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__5180__A1 _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5823__I _4529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8957__B1 _3993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5698__C _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8421__A2 _3361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5235__A2 _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8488__A2 _3366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6499__A1 _4541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5171__A1 _4518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5733__I _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8660__A2 _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5474__A2 _4478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6564__I _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6423__A1 as2650.stack\[2\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5401__C _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5971_ _1234_ _1236_ _1244_ _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_52_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7710_ as2650.pc\[7\] net2 _2842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4922_ _4356_ _4502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8690_ _1624_ _4377_ _3778_ _1535_ _3779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__8176__A1 _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7641_ _2520_ _2774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4853_ _4426_ _4433_ _4434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7395__I _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7923__A1 _3048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6726__A2 _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7572_ _0507_ _0490_ _2671_ _2672_ _2707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__9166__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4784_ _4320_ _4365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_18_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9311_ _0204_ clknet_3_3_0_wb_clk_i as2650.cycle\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
X_6523_ _1750_ _1755_ _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_140_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8479__A2 _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9242_ _0135_ clknet_leaf_55_wb_clk_i as2650.stack\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6454_ _1239_ _1690_ _1694_ _0071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7151__A2 _2248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5405_ _0711_ _0343_ _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5162__A1 _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9173_ _0066_ clknet_leaf_60_wb_clk_i as2650.stack\[2\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6385_ _0851_ _1640_ _1019_ _1641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_8124_ _3230_ _3231_ _3233_ _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5336_ _0567_ _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_142_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8100__A1 _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8055_ _3158_ _1370_ _3159_ _3167_ _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__8651__A2 _3727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5267_ _0290_ _0481_ _0502_ _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_29_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7006_ _2204_ _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5799__B _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5198_ _0506_ _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6474__I _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6414__A1 _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8957_ _0703_ _3992_ _3993_ as2650.r123\[2\]\[5\] _4002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7908_ as2650.pc\[12\] _3035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_24_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8888_ as2650.stack\[7\]\[9\] _3951_ _3952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8622__C _3048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7839_ _0988_ _2968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_70_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7914__A1 _3018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4728__A1 _4291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7390__A2 _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5153__A1 _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6350__B1 _4526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5553__I _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6350__C2 _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8642__A2 _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6248__A4 _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6384__I _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5208__A2 _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5759__A3 _4245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6956__A2 _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9189__CLK clknet_leaf_65_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5392__A1 _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8330__A1 _3428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6341__B1 _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6170_ _0569_ _0662_ _0740_ _1427_ _1428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_124_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5121_ as2650.stack\[0\]\[10\] _0429_ _0430_ as2650.stack\[1\]\[10\] _0431_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_123_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6495__I1 as2650.r123_2\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7611__C _2744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5052_ as2650.r0\[3\] _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4807__I _4387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6294__I _4531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8811_ _2109_ _3844_ _3847_ _3892_ _1624_ _3893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_93_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8742_ as2650.psu\[3\] _3771_ _3828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5954_ _1227_ _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8149__A1 _3208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4905_ _4472_ _4484_ _4485_ _4486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8673_ _3219_ _4344_ _3183_ _3760_ _3761_ _3762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5885_ _4228_ _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5638__I _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7624_ _2757_ _2504_ _2688_ _2736_ _2529_ _2758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4836_ _4170_ _4417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7372__A2 _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7555_ _2689_ _2649_ _2690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4767_ _4243_ _4347_ _4348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6506_ _1739_ _1740_ _0077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7486_ _2529_ _2617_ _2622_ _2623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8321__A1 _2416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7124__A2 _2286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4698_ _4277_ _4278_ _4279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5135__A1 _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9225_ _0118_ clknet_leaf_55_wb_clk_i as2650.stack\[4\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6437_ _1335_ _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5373__I _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9156_ _0049_ clknet_leaf_56_wb_clk_i as2650.stack\[4\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6368_ _1622_ _1624_ _1625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8107_ _3211_ _3213_ _3215_ _3216_ _3217_ _3218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_62_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5319_ as2650.stack\[0\]\[12\] _4482_ _0626_ as2650.stack\[1\]\[12\] _0627_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_49_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9087_ _4108_ _4117_ _4118_ _3249_ _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_114_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6299_ _1551_ _1552_ _1555_ _1556_ _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_130_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5438__A2 _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8038_ _3106_ _3151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9331__CLK clknet_leaf_80_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6932__I _4295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5548__I _4204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8560__A1 _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8859__I _3926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8312__A1 _3070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8795__S _3792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5429__A2 _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4627__I as2650.cycle\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8379__A1 _3459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5659__S _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8035__S _3119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5670_ _0965_ _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8551__A1 _2969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7354__A2 _4393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4621_ net5 _4202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7340_ _1678_ _1676_ _4240_ _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_11_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5407__B _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7271_ _1356_ _1513_ _2410_ _1370_ _2411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__9204__CLK clknet_leaf_46_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9010_ _3214_ _1551_ _3126_ _1249_ _4048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_137_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6222_ _1044_ _1480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_144_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5912__I0 _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_49_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6153_ _1416_ _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6617__A1 as2650.r0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9354__CLK clknet_leaf_59_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5104_ _0314_ _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6084_ _1355_ _1305_ _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6238__B _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7290__A1 _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5035_ _4500_ _0323_ _0345_ _4498_ _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_100_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9031__A2 _3074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7042__A1 _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6986_ _2187_ _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8790__A1 _3837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5937_ _0473_ _0801_ _1210_ _1211_ _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
X_8725_ as2650.overflow _3812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_107_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8656_ _2755_ _0600_ _3744_ _3175_ _4260_ _3745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_5868_ _0508_ _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8542__A1 _3625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7607_ _2706_ _2739_ _2707_ _2740_ _2741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_55_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4819_ _4398_ _4399_ _4400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8587_ _3153_ _3672_ _3679_ _3680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6553__B1 _1784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5799_ _4353_ _1057_ _1080_ _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7538_ _1585_ _0491_ _2673_ _2674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_33_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4954__I1 _4533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7469_ _2602_ _2605_ _2606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_134_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput13 net50 io_oeb[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__6856__A1 _4367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput24 net24 io_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_9208_ _0101_ clknet_leaf_77_wb_clk_i as2650.r123_2\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput35 net35 io_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__4706__I1 as2650.r123\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9139_ _0032_ clknet_leaf_46_wb_clk_i as2650.r123_2\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8347__C _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6084__A2 _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7281__A1 _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7820__A3 _2869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9022__A2 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7033__A1 _2183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8781__A1 _3769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8781__B2 _3847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5595__A1 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5595__B2 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5278__I _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7493__I _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4910__I _4490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5898__A2 _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9089__A2 _2925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4570__A2 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8836__A2 _3912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6847__A1 _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9377__CLK clknet_leaf_9_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7272__A1 _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9013__A2 _3113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6840_ _2021_ _2047_ _2050_ _2051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_63_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7575__A2 _2585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8772__A1 _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5586__A1 _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6771_ _1944_ _1978_ _1983_ _1984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_50_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8510_ _3533_ _3602_ _3604_ _3605_ _3606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_17_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4928__A4 _4385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5722_ as2650.stack\[6\]\[13\] _0962_ _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_31_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8441_ _2800_ _0583_ _3539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5653_ _0950_ _0014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5916__I as2650.r123_2\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4604_ _4181_ _4184_ _4185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_8372_ _2648_ _3469_ _3470_ _3471_ _3472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5584_ _4251_ _4164_ _0884_ _0887_ _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_141_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7323_ _2437_ _2438_ _2461_ _2462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_89_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_5_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6838__A1 _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7254_ _2395_ _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6302__A3 _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6205_ _1462_ _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7185_ _1272_ _2335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6136_ _1399_ _0593_ _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6066__A2 _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8460__B1 _3557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6067_ _0881_ _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5813__A2 _4261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5018_ _0328_ _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7015__A1 _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8763__A1 _3844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8763__B2 _3847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6969_ _2170_ _2171_ _2172_ as2650.stack\[2\]\[1\] _2173_ _2174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_41_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8708_ _1733_ _3769_ _4435_ _3795_ _3777_ _3796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_70_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8515__A1 _2899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7318__A2 _4443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8639_ _1008_ _3707_ _3729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8818__A2 _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5501__A1 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5561__I _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6057__A2 _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8093__B _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5510__B _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5280__A3 _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7557__A2 _2688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8754__A1 _3804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5568__A1 _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8506__A1 _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7309__A2 _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7951__I _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8809__A2 _3793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4796__B _4321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input1_I io_in[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6048__A2 _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8990_ _0854_ _4030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8993__A1 _4010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7941_ _4169_ _2348_ _3066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7398__I _4531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7260__A4 _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7872_ _2995_ _2996_ _2997_ _2999_ _3000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_70_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8745__A1 _3826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6823_ _0362_ _1965_ _2035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8731__B _3817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6220__A2 _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6754_ _1842_ _1966_ _1967_ _1881_ _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__8450__C _3154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5705_ _0441_ _0981_ _0982_ _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6685_ as2650.stack\[1\]\[9\] _1911_ _1912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5646__I _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8424_ as2650.stack\[4\]\[5\] _1904_ _1656_ as2650.stack\[5\]\[5\] _3523_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_5636_ _0915_ _0935_ _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8355_ _0927_ _3423_ _3455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5567_ _0870_ _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7306_ _2436_ _2441_ _2442_ _2444_ _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_132_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8286_ _0327_ _3387_ _3388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5498_ _0724_ _0794_ _0797_ _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7237_ _1309_ _1491_ _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6477__I _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7168_ _2258_ _2318_ _2319_ as2650.stack\[0\]\[2\] _2320_ _2324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_144_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7236__A1 _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6039__A2 _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6119_ _4202_ _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7099_ as2650.r123\[3\]\[2\] _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8625__C _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8984__A1 _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5798__A1 _4361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7539__A2 _2674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8736__A1 _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6211__A2 _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6940__I _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5970__A1 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5556__I _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7711__A2 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5722__A1 as2650.stack\[6\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8088__B _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6278__A2 _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8816__B _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8424__B1 _1656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7778__A2 _2684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8727__A1 _3812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6202__A2 _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7950__A2 _3074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6470_ _1707_ _0074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7702__A2 _2704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5421_ _0642_ _0644_ _0659_ _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5713__A1 _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5713__B2 as2650.r123_2\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8140_ as2650.cycle\[5\] _3247_ _3248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_103_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5352_ _0637_ _0638_ _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6297__I _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8071_ _3183_ _3184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5283_ _0590_ _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_134_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7022_ _2213_ _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7769__A2 _2532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8966__A1 _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8445__C _3070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8973_ _2409_ _1481_ _4013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6441__A2 _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7924_ _1331_ _2412_ _3047_ _3049_ _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_70_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7855_ _2945_ _2946_ _2983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8194__A2 _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6806_ _1982_ _2018_ _0099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7786_ _2361_ _2879_ _2916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5401__B1 _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4998_ _4315_ _0308_ _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7941__A2 _2348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6737_ _1879_ _1885_ _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5376__I _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6668_ _1867_ _1896_ _1897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_104_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8351__C1 _3451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5619_ _0920_ _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8407_ _2694_ _0496_ _3506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_118_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6599_ _1782_ _1802_ _1829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9387_ _0280_ clknet_leaf_5_wb_clk_i as2650.psl\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8338_ _3400_ _3404_ _3438_ _3439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7457__A1 _4528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8269_ _3337_ _3370_ _3371_ _3372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_79_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4691__A1 _4154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8957__A1 _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output40_I net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6432__A2 _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8709__A1 _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6196__A1 _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5943__A1 _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4746__A2 _4325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5286__I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7696__A1 _1617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6499__A2 _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5171__A2 _4523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_57_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_57_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_124_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7006__I _2204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6671__A2 _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4682__A1 _4235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8412__A3 _3428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5970_ _1237_ _1241_ _1243_ _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_93_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4921_ _4408_ _4501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8281__B _4473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8176__A2 _2506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7640_ _2579_ _2770_ _2773_ _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_33_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6187__A1 _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4852_ _4427_ _4430_ _4432_ _4433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__9096__C _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7923__A2 _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7571_ _0507_ _0490_ _2706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4783_ _4221_ _4364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5934__A1 _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5196__I _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4737__A2 _4311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9310_ _0203_ clknet_leaf_18_wb_clk_i as2650.cycle\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6522_ _0364_ _1722_ _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7687__A1 _2751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9241_ _0134_ clknet_leaf_55_wb_clk_i as2650.stack\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6453_ _1552_ _1692_ _1689_ _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5404_ _0670_ _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_9172_ _0065_ clknet_leaf_60_wb_clk_i as2650.stack\[2\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5162__A2 _4422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6384_ _1639_ _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8123_ _0893_ _3232_ _3233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_114_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5335_ as2650.holding_reg\[5\] _0591_ _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_138_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8100__A2 _3090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8054_ _1676_ _1236_ _1249_ _3166_ _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_134_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5266_ _0290_ _0481_ _0502_ _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_7005_ _2203_ _2204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6662__A2 _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5197_ net9 _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4673__A1 _4163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7611__A1 _2704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8956_ _3976_ _2100_ _4001_ _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7907_ _2923_ _3029_ _3033_ _3034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_8887_ _3946_ _3951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8167__A2 _3271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6178__A1 _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7838_ _2923_ _2966_ _2967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_58_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9110__CLK clknet_leaf_68_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5925__A1 _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4728__A2 _4256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7769_ _2884_ _2532_ _2535_ _2899_ _2502_ _2900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_32_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9260__CLK clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6350__A1 _4530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5153__A2 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6350__B2 _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8627__B1 _3712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6102__A1 _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5759__A4 _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7496__I _2631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6169__A1 _4344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8563__C1 _3103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5392__A2 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7445__B _2581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8330__A2 _3429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8120__I _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7164__C _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5144__A2 _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6341__A1 as2650.psl\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6341__B2 _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6892__A2 _1942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_39_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5120_ _4469_ _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8094__A1 _3201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7841__A1 _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5051_ _0360_ _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8810_ _3262_ _3793_ _3891_ _3892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_92_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8741_ _4365_ _3827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_92_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5953_ _0876_ _4157_ _4278_ _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5080__A1 _4354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8149__A2 _2484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4904_ _4445_ _4485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5884_ _0603_ _1070_ _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8672_ _3143_ _1100_ _3080_ _3761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_94_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7623_ net33 _2757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__9283__CLK clknet_leaf_26_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4835_ _4415_ _4416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5907__A1 _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7554_ net31 _2689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4766_ as2650.idx_ctrl\[0\] _4347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_140_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6505_ _1116_ _1717_ _1740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7485_ _2609_ _2618_ _2500_ _2621_ _2622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_119_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4697_ _4159_ _4178_ _4278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5654__I _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8321__A2 _3422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9224_ _0117_ clknet_leaf_39_wb_clk_i as2650.stack\[4\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7074__C _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6436_ _1464_ _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_9155_ _0048_ clknet_leaf_57_wb_clk_i as2650.stack\[4\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6367_ _1623_ _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4894__A1 _4473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8106_ _3211_ _3213_ _3217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8085__A1 _3164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5318_ _0324_ _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6298_ _1147_ _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_9086_ _4041_ _4108_ as2650.psl\[1\] _4118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6485__I _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6635__A2 _1858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8037_ _2416_ _1488_ _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5249_ _0444_ _0453_ _0466_ _0442_ _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_5_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4646__A1 _4181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_2_wb_clk_i clknet_3_0_0_wb_clk_i clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_29_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6399__A1 _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8939_ _3988_ _3989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5071__A1 _4378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4733__I _4313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7899__A1 _2662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7899__B2 _2476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8560__A2 _2776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6571__A1 _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5564__I _4215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8312__A2 _3407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5126__A2 _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7823__A1 _2866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6626__A2 _1849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9156__CLK clknet_leaf_56_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7587__B1 _2718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8543__C _2928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8115__I _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8551__A2 _3644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4620_ _4200_ _4201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_2
XFILLER_19_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6562__A1 _1174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7270_ _0896_ _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_132_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6221_ _1465_ _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_116_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8067__A1 _3178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6152_ _1416_ _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5103_ as2650.holding_reg\[2\] _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7814__A1 _2919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6617__A2 _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4818__I _4396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6083_ _1355_ _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5034_ _4494_ _0336_ _0344_ _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_39_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7290__A2 _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9031__A3 _4067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7042__A2 _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6985_ as2650.pc\[4\] _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5649__I _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4553__I net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8790__A2 _3872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8724_ _0618_ _3390_ _3811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5936_ _0473_ _0819_ _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8655_ _1329_ _2472_ _3265_ _3744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5867_ _4188_ _1040_ _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__8542__A2 _3627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7606_ _0595_ _0577_ _2740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4818_ _4396_ _4399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8586_ _3674_ _3677_ _3678_ _3679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5798_ _4361_ _1059_ _1060_ _1079_ _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_120_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7537_ _2671_ _2672_ _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4749_ _4329_ _4330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6305__A1 _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7468_ _2568_ _2603_ _2604_ _2605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput14 net14 io_oeb[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_9207_ _0100_ clknet_leaf_77_wb_clk_i as2650.r123_2\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput25 net25 io_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__6856__A2 _1764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6419_ _0992_ _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput36 net36 io_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_7399_ _2530_ _2417_ _2537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_66_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9179__CLK clknet_leaf_9_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8058__A1 _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9138_ _0031_ clknet_leaf_46_wb_clk_i as2650.r123_2\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6608__A2 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9069_ _2793_ _1469_ _4103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7281__A2 _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6943__I _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7033__A2 _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5559__I _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9178__D _0071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8781__A2 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5595__A2 _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6544__A1 _1757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8297__A1 _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6847__A2 _2027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8049__A1 _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7014__I _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7272__A2 _2408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7949__I _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8221__A1 as2650.stack\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8772__A2 _3856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5586__A2 _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6770_ _1945_ _1946_ _1977_ _1983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5721_ _1011_ _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_91_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8440_ _2800_ _0583_ _3538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6535__A1 _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5652_ _0944_ _0949_ _0860_ _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_30_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4603_ _4155_ _4183_ _4184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5583_ _4234_ _0885_ _0886_ _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_8371_ _1267_ _0898_ _3471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7322_ _4161_ _2458_ _0833_ _2460_ _2461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__9321__CLK clknet_leaf_31_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6838__A2 _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7253_ _4176_ _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6204_ _4250_ _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7184_ _2333_ _2334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5510__A2 _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6135_ _1397_ _1401_ _1403_ _1392_ _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_131_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6066_ _1336_ _1338_ _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8460__A1 _3216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8460__B2 _3481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5274__A1 _4521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5017_ _0327_ _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8212__A1 _3214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8763__A2 _2027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6968_ _2141_ _2173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8707_ _4458_ _3793_ _3794_ _3795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5919_ _0753_ _1103_ _1066_ _1194_ _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6899_ _2106_ _2107_ _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8515__A2 _3610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7318__A3 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8638_ _4264_ _3158_ _3625_ _3728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_139_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8569_ _2969_ _3621_ _3662_ _3592_ _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_33_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8279__A1 _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6003__I _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6938__I _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7262__C _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5501__A2 _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8451__A1 _3153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5265__A1 _4359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8203__A1 _4161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5289__I _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8754__A2 _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5568__A2 _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6765__A1 _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8506__A2 _2903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7309__A3 _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4921__I _4408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9344__CLK clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5740__A2 _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5752__I _4200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8690__A1 _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8993__A2 _4028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7940_ _1356_ _1684_ _1504_ _3065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_36_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7871_ _2982_ _2504_ _2507_ _2998_ _1268_ _2999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_58_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5199__I _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5008__A1 _4338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6822_ _2004_ _2008_ _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8731__C _3765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6753_ _1880_ _1883_ _1967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_50_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4831__I _4262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5704_ _0996_ _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6508__A1 _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6684_ _1906_ _1911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8423_ as2650.stack\[7\]\[5\] _3366_ _3386_ as2650.stack\[6\]\[5\] _3522_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_5635_ _0933_ _0903_ _0934_ _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7181__A1 _2307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8354_ _0928_ _3289_ _3454_ _3112_ _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_30_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5731__A2 _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5566_ _4255_ _0869_ _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7305_ _1346_ _1683_ _2443_ _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_105_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9281__D _0174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5497_ _0796_ _0798_ _0801_ _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8285_ as2650.stack\[7\]\[2\] _1918_ _1902_ as2650.stack\[4\]\[2\] as2650.stack\[5\]\[2\]
+ _1654_ _3387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_104_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7484__A2 _2620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7236_ _2377_ _2358_ _2378_ _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8681__A1 _4428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7082__C _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7167_ _2321_ _2323_ _0155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_28_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6118_ net43 _1380_ _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8433__A1 _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7236__A2 _2358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6039__A3 _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7098_ _2270_ _0139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8984__A2 _4020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6049_ _1315_ _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5798__A2 _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8736__A2 _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9367__CLK clknet_leaf_68_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4758__B1 _4336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8213__I _2387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7257__C _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5970__A2 _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7172__A1 _2298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5722__A2 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7273__B _2412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5572__I _4180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8088__C _3199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8672__A1 _3143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8883__I _3947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8424__B2 as2650.stack\[5\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7499__I _2634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8727__A2 _3772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7448__B _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5410__A1 _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7950__A3 _2412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5420_ _0555_ _0724_ _0725_ _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_127_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6910__A1 _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5351_ _0646_ _0650_ _0657_ _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_142_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8112__B1 _2508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5482__I _4494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7466__A2 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8663__A1 _4242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8070_ _3182_ _3183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5282_ _0589_ _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_47_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5477__A1 _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7021_ _2138_ _2211_ _2218_ _0114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_87_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8415__A1 _3059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8966__A2 _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8972_ _2926_ _4011_ _4012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout52_I net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7923_ _3048_ _2152_ _4444_ _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_97_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8718__A2 _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7854_ net39 _2982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8461__C _3288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6805_ _1727_ _2017_ _2018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7785_ _2912_ _2914_ _2915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_24_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5401__A1 as2650.stack\[3\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4997_ _0305_ _0307_ _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5401__B2 as2650.stack\[2\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6736_ _1879_ _1885_ _1950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6667_ _1870_ _1895_ _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_137_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8351__C2 _3327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8406_ _2694_ _0496_ _3505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5618_ _0919_ _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6901__A1 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9386_ _0279_ clknet_leaf_3_wb_clk_i as2650.psl\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_87_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6598_ _1785_ _1786_ _1828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8337_ _3399_ _3438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5549_ _4487_ _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7457__A2 _4511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8654__A1 _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8268_ _3290_ _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5468__A1 _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7219_ _2366_ _2363_ _2367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4937__S _4516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8199_ _2458_ _0834_ _2460_ _3303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_8_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8406__A1 _2694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7540__C _2564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8957__A2 _3992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4691__A2 _4189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7112__I _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output33_I net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8709__A2 _4514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6951__I _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6196__A2 _4541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7393__A1 _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5567__I _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5943__A2 _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7145__A1 _2200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7696__A2 _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8893__A1 _1668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_29_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5171__A3 _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_3_6_0_wb_clk_i clknet_0_wb_clk_i clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_123_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5459__A1 _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_0_wb_clk_i_I wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_26_wb_clk_i clknet_opt_1_0_wb_clk_i clknet_leaf_26_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__9070__A1 _3770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8118__I _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7022__I _2213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7957__I _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4920_ _4274_ _4500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4851_ _4312_ _4431_ _4432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_127_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7570_ _2565_ _2704_ _2705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4782_ _4362_ _4363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_68_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6521_ _1139_ _1715_ _1754_ _0078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7136__A1 _2298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9240_ _0133_ clknet_leaf_38_wb_clk_i as2650.stack\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7687__A2 _2813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6452_ _1523_ _1690_ _1693_ _0070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5698__A1 _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5698__B2 as2650.r123_2\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5403_ _4485_ _0709_ _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_9171_ _0064_ clknet_leaf_60_wb_clk_i as2650.stack\[2\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6383_ _1638_ _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6101__I _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8122_ _3209_ _1507_ _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8636__A1 _3724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5334_ _0640_ _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8053_ _1237_ _1045_ _1273_ _3166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_87_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5265_ _4359_ _0503_ _0573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_102_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7004_ as2650.pc\[7\] _2203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5196_ _0504_ _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4673__A2 _4253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5870__A1 _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8028__I _3143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9061__A1 _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7611__A2 _2742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8955_ _0616_ _3986_ _3989_ as2650.r123\[2\]\[4\] _4001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8472__B _3504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7867__I _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7906_ _2607_ _3032_ _3033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8886_ _1653_ _3948_ _3950_ _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7837_ _2658_ _2964_ _2965_ _2966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_24_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5387__I _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7768_ _2866_ _2899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_71_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6719_ _1674_ _1925_ _1933_ _0097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7127__A1 _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7699_ _0757_ _0771_ _2831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9438_ net46 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8875__A1 _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5689__A1 _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5689__B2 as2650.r123_2\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9369_ _0262_ clknet_leaf_74_wb_clk_i as2650.r123\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_4_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6350__A2 _4387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8627__A1 _3257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8627__B2 _2549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7850__A2 _2967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9052__A1 _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8382__B _4473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6681__I _1907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6169__A2 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7118__A1 _2147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8315__B1 _3414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7118__B2 as2650.stack\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8866__A1 _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6341__A2 _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7017__I _4474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5050_ _0359_ _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7180__C _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4655__A2 as2650.cycle\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5852__A1 _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5604__A1 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8740_ _0618_ _3451_ _3826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_81_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5952_ as2650.psu\[5\] _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5080__A2 _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4903_ _4477_ _4480_ _4483_ _4484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_8671_ _2477_ _4353_ _3759_ _3760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7357__A1 _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5883_ _0617_ _0621_ _0632_ _1088_ _1090_ _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_59_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7622_ _2755_ _2756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4834_ _4205_ _4415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7553_ _2507_ _2688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4765_ _4345_ _4346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6504_ as2650.r123_2\[1\]\[1\] _1729_ _1727_ _1738_ _1739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_135_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8857__A1 _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7484_ _1545_ _2620_ _2621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8857__B2 as2650.stack\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4696_ _4192_ _4277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9223_ _0116_ clknet_leaf_40_wb_clk_i as2650.stack\[4\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6435_ _1676_ _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_134_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8609__A1 _3210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9154_ _0047_ clknet_leaf_57_wb_clk_i as2650.stack\[4\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6366_ _4219_ _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8105_ _2388_ _3216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4894__A2 _4474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6766__I _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5317_ as2650.stack\[2\]\[12\] _0624_ _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9085_ _1382_ _4113_ _4116_ _4117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6297_ _1554_ _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6096__A1 _4328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8036_ _3150_ _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7090__C _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5248_ _0549_ _0504_ _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_88_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9034__A1 _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5179_ _0477_ _0478_ _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7596__A1 _2728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8938_ _1390_ _3961_ _3985_ _3988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_45_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5071__A2 _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7348__A1 _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8869_ _2296_ _3931_ _3932_ as2650.stack\[7\]\[3\] _3933_ _3939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_52_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8848__A1 _2307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7520__A1 _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5580__I as2650.cycle\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6087__A1 _4215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7823__A2 as2650.addr_buff\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5834__A1 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9025__A1 _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7036__B1 _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7587__A1 _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7587__B2 _2719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7339__A1 _2467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7339__B2 _2477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6011__A1 _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7456__B _4528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6562__A2 _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4573__A1 _4143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8839__A1 _2298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7511__A1 _2643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7970__I _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6220_ _4187_ _1477_ _4419_ _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7191__B _1496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6151_ _1415_ _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_41_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_41_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5490__I _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6078__A1 _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5102_ _0409_ _0410_ _0411_ _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_98_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7814__A2 _2942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6082_ _4207_ _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4628__A2 _4208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5825__A1 _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5033_ _0337_ _0343_ _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_61_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9016__A1 _3492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6984_ _0617_ _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6250__A1 _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8723_ _1623_ _3810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5935_ _1208_ _1209_ _0815_ _0651_ _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_22_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4800__A2 _4380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8654_ _1453_ _2420_ _3743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5866_ _1082_ _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_61_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7605_ _0595_ _0577_ _2739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_107_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4817_ _4216_ _4333_ _4398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8585_ _3256_ _3664_ _3673_ _2524_ _2927_ _3678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_33_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7750__A1 _2334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5797_ _1061_ _1078_ _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8041__I _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7536_ _0374_ _2592_ _2593_ _2561_ _2594_ _2672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_4748_ _4323_ _4328_ _4329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7467_ _0909_ net7 _2604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7502__A1 _2636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4679_ _4254_ _4259_ _4260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_123_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9206_ _0099_ clknet_leaf_73_wb_clk_i as2650.r123_2\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_123_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6418_ _1663_ _1660_ _1665_ _0064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xoutput15 net15 io_oeb[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_135_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput26 net26 io_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_7398_ _4531_ _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput37 net37 io_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__4706__I3 as2650.r123_2\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6496__I _1730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9137_ _0030_ clknet_leaf_46_wb_clk_i as2650.r123_2\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6349_ _1549_ _4334_ _0592_ _0684_ _0753_ _1605_ _1606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_88_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6069__A1 _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9068_ _3812_ _4097_ _4102_ _3249_ _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_131_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9007__A1 _3230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8019_ _1558_ _3136_ _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7281__A3 _2419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8216__I _1654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7120__I _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6241__A1 _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8660__B _4395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5595__A3 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7741__A1 _2871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5575__I _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6544__A2 _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8297__A2 _4517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9123__CLK clknet_leaf_58_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8049__A2 _2348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9273__CLK clknet_leaf_12_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6480__A1 _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8757__B1 _3184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8221__A2 _3322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5035__A2 _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_63_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7965__I _3089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7980__A1 _3103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5720_ _1008_ _0858_ _0972_ as2650.r123_2\[0\]\[5\] _1010_ _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_108_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5651_ _0948_ as2650.stack\[5\]\[6\] _0902_ _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5485__I _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7732__A1 _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4602_ _4182_ _4183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8370_ _0596_ _1490_ _3470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5582_ _4239_ _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_129_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7321_ _0512_ _0603_ _0690_ _2459_ _2460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_102_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6299__A1 _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7252_ _1366_ _2379_ _2393_ _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_116_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6203_ _1451_ _1460_ _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7183_ as2650.addr_buff\[0\] _2333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6134_ net45 _1402_ _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7799__A1 _2777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8745__B _3777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6065_ _4238_ _1337_ _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5274__A2 _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5016_ _4453_ _4451_ _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__9279__D _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4564__I _4144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6223__A1 _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6967_ _2167_ _2172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7971__A1 net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5918_ _0759_ _1105_ _1193_ _1165_ _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_8706_ as2650.psl\[1\] _3792_ _3794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6898_ _2079_ _2089_ _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7318__A4 _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8637_ _3726_ _3727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5849_ _0376_ _1105_ _1128_ _1102_ _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7723__A1 _1497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8920__B1 _3964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9146__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8568_ _3379_ _3645_ _3660_ _3661_ _3373_ _3662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7519_ _2335_ _2527_ _2655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7824__B _2564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8499_ _0965_ _3594_ _3595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_68_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7543__C _2483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4739__I as2650.psl\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7115__I _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8655__B _3265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6954__I _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5265__A2 _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7962__A1 _2463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7309__A4 _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7714__A1 _2837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7714__B2 _2818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8911__B1 _3967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5725__B1 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8549__C _3592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4649__I _4229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8690__A2 _4377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6453__A1 _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7870_ as2650.addr_buff\[3\] _2998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_36_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6821_ _2031_ _2032_ _2033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7953__A1 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6752_ as2650.r0\[1\] _1965_ _1966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9169__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5703_ _0995_ _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_91_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6683_ _1653_ _1908_ _1910_ _0084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_32_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8422_ _3518_ _0426_ _3519_ _4453_ _3520_ _3521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__6104__I _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5634_ as2650.stack\[5\]\[4\] _0913_ _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8353_ _3333_ _3425_ _3453_ _3454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5192__A1 _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5565_ _4224_ _4369_ _4313_ _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_129_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7304_ _1497_ _4250_ _2443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8284_ _1637_ _3386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8130__A1 _2624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5496_ _0800_ _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_104_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7235_ _1340_ _2363_ _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_137_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6692__A1 _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5495__A2 _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7166_ _2290_ _2322_ _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8475__B _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6117_ _0917_ _1376_ _1387_ _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8433__A2 _1618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7097_ as2650.r123\[3\]\[1\] _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6444__A1 _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6048_ _1320_ _1228_ _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_86_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8984__A3 _4022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8197__A1 as2650.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7944__A1 _2349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6747__A2 _1730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6723__B _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7999_ _3115_ _4291_ _3120_ _3121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_96_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4758__A1 _4330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5970__A3 _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6014__I _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7273__C _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8121__A1 _1681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8672__A2 _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6683__A1 _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8424__A2 _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9311__CLK clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_58_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7950__A4 _2451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5174__A1 _4524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5350_ _0651_ _0653_ _0656_ _0553_ _0562_ _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__8112__A1 _4253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8112__B2 _3059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8663__A2 _2469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5281_ _0588_ _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_141_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7020_ _2147_ _2214_ _2217_ as2650.stack\[4\]\[0\] _2210_ _2218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__7871__B1 _2507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6426__A1 as2650.stack\[2\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8971_ _3191_ _2509_ _3048_ _1309_ _4011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_82_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7922_ _0871_ _3048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4988__A1 _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8179__A1 _4444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7853_ _2521_ _2980_ _2981_ _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_82_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6729__A2 _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6804_ _1984_ _2016_ _2017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_24_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7784_ _2913_ _2895_ _2914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4996_ _4317_ _0306_ _4310_ _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5401__A2 _4479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6735_ _1888_ _1892_ _1948_ _1949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6666_ _1873_ _1894_ _1895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8351__A1 _3426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7154__A2 _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8351__B2 _3446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5617_ as2650.pc\[2\] _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8405_ _3471_ _3504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5165__A1 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9385_ _0278_ clknet_leaf_71_wb_clk_i as2650.psl\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6597_ _1798_ _1822_ _1826_ _1827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5673__I _4152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6901__A2 _2109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8336_ _3156_ _3425_ _3431_ _3436_ _3437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4912__A1 _4415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5548_ _4204_ _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_133_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8267_ _3199_ _3359_ _3368_ _3369_ _3370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7457__A3 _4512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5479_ _4274_ _0775_ _0784_ _0538_ _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_69_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8654__A2 _2420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5468__A2 _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7218_ _2365_ _2366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8198_ _3296_ _3301_ _3302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_115_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8406__A2 _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7149_ _2307_ _2291_ _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9334__CLK clknet_leaf_80_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7090__A1 _2265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6009__I _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output26_I net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7917__A1 _2521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4752__I _4304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8590__A1 _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6196__A3 _4405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout50 net13 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_70_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8342__A1 _2854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8893__A2 _3948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_6_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4903__A1 _4477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5171__A4 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4927__I _4506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4682__A3 _4240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9070__A2 _3268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_66_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_66_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_3392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7178__C _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4850_ _4156_ _4313_ _4431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_60_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8581__A1 _3533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6187__A3 _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5395__A1 _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4781_ _4213_ _4362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6520_ as2650.r123_2\[1\]\[2\] _1719_ _1741_ _1753_ _1754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_18_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8333__A1 _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7136__A2 _2291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9207__CLK clknet_leaf_77_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6451_ _1691_ _1692_ _1690_ _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5402_ _0704_ _0705_ _0708_ _0526_ _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_134_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9170_ _0063_ clknet_leaf_60_wb_clk_i as2650.stack\[2\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6382_ _1637_ _1638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8121_ _1681_ _2155_ _3221_ _3231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5333_ _0637_ _0639_ _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_86_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8737__C _2756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6647__A1 as2650.r0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8052_ _2535_ _3162_ _3164_ _3165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__9357__CLK clknet_leaf_60_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5264_ _0477_ _0541_ _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_69_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7003_ _2200_ _2143_ _2202_ _0112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4837__I _4417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7213__I _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5195_ _0503_ _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_60_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5870__A2 _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9061__A2 _4010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8954_ _3999_ _4000_ _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8472__C _3568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7905_ _3012_ _3031_ _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_97_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5668__I as2650.pc\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8885_ as2650.stack\[7\]\[8\] _3949_ _3950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8044__I _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7836_ _2962_ _2963_ _2960_ _2965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7767_ _2895_ _2897_ _2751_ _2898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4979_ _4508_ _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6718_ as2650.stack\[0\]\[14\] _1923_ _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_71_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7698_ _2588_ _2828_ _2829_ _2554_ _2830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7127__A2 _2291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9437_ net47 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6649_ _1876_ _1877_ _1878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6335__B1 _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9368_ _0261_ clknet_leaf_65_wb_clk_i as2650.r123\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7832__B _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8319_ _3379_ _3418_ _3419_ _3420_ _3421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_133_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8627__A2 _3706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9299_ _0192_ clknet_leaf_1_wb_clk_i as2650.holding_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_59_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8647__C _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7123__I _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8663__B _3751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6962__I _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5578__I _4254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8563__A1 _3504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6169__A3 _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8563__B2 _3459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7793__I _2570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8315__A1 _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8315__B2 _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6326__B1 _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8866__A2 _3931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6877__A1 _4367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7968__I _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5951_ _1205_ _1160_ _1225_ _0037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4902_ as2650.stack\[4\]\[8\] _4482_ _4470_ as2650.stack\[5\]\[8\] _4483_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8670_ _2598_ _4361_ _3759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5882_ _1054_ _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7357__A2 _2495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7621_ _2754_ _2755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4833_ _4276_ _4344_ _4413_ _4414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__5368__A1 _4369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7552_ net32 _2687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4764_ _4247_ _4345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8306__A1 _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6503_ _1735_ _1737_ _1738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7483_ _2602_ _2619_ _2620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_119_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4695_ _4262_ _4276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_135_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7208__I _2357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6434_ _1500_ _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_9222_ _0115_ clknet_leaf_40_wb_clk_i as2650.stack\[4\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8748__B _2629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9153_ _0046_ clknet_leaf_16_wb_clk_i net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8609__A2 _3686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6365_ _1442_ _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5540__A1 _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8104_ _1304_ _4175_ _3214_ _3215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5316_ _4460_ _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_66_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9084_ _1552_ _3136_ _4100_ _4116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_130_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6296_ _1553_ _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_27_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4567__I _4147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8035_ _3149_ _0813_ _3119_ _3150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6096__A2 _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5247_ _4315_ _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4646__A3 _4226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9034__A2 _4056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5178_ _4359_ _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_60_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7596__A2 _2729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8793__A1 _2635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8937_ _3986_ _3987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_44_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8868_ _3937_ _3938_ _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7348__A2 _4391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7827__B _2366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5359__A1 _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7819_ _2744_ _2876_ _2878_ _2948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_8799_ _3767_ _0818_ _3780_ _3882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_40_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8848__A2 _3912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7520__A2 _2655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7284__A1 _4427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5834__A2 _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9025__A2 _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8393__B _3288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7036__A1 _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7587__A2 _2715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5047__B1 _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8784__A1 _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5598__A1 _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8536__A1 _3221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7737__B _4245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4940__I _4519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4573__A2 _4153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8839__A2 _3912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7511__A2 _2644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6150_ _0622_ _1019_ _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_139_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6078__A2 _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5101_ _4277_ _4324_ _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_83_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6081_ _4168_ _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5032_ _0342_ _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5825__A2 _4534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9016__A2 _4051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7027__A1 _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8224__B1 _3326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7578__A2 _2712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8775__A1 _3804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6983_ _2184_ _2185_ _0109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6250__A2 _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6107__I _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8722_ _0378_ _2632_ _3809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5934_ _0544_ _0807_ _0812_ _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8653_ _3724_ _3621_ _3741_ _3742_ _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5865_ _0536_ _1117_ _1143_ _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_90_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7604_ _2588_ _2735_ _2737_ _2662_ _2738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4816_ _4396_ _4397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8584_ _2495_ _3665_ _3675_ _1277_ _3676_ _3677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_22_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5796_ _4406_ _1063_ _1077_ _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7535_ _0375_ _2592_ _2671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4747_ _4178_ _4328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5761__A1 _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7466_ as2650.pc\[1\] net7 _2603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4678_ _4198_ _4257_ _4245_ _4258_ _4259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6417_ as2650.stack\[2\]\[9\] _1664_ _1665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_9205_ _0098_ clknet_leaf_74_wb_clk_i as2650.r123_2\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7397_ _2534_ _2535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5681__I _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput16 net16 io_oeb[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput27 net27 io_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_1_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput38 net38 io_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_6348_ _1604_ _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_9136_ _0029_ clknet_leaf_58_wb_clk_i as2650.stack\[5\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9067_ _4098_ _4099_ _4101_ _1576_ _4097_ _4102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_6279_ _0718_ _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8018_ _2794_ _3136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_44_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9007__A2 _4040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7018__A1 _2215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7401__I _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6241__A2 _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6017__I _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8518__A1 _3257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8518__B2 _2550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5856__I _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7741__A2 _2869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7292__B _2406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8835__C _3910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6480__A2 _4489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8757__A1 _3838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8509__A1 _2996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_50_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7980__A2 _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5991__A1 _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9385__D _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4670__I as2650.cycle\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8142__I _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5650_ _0947_ _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7732__A2 _2580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4601_ as2650.ins_reg\[5\] _4182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5581_ _4238_ _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5743__A1 _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7320_ _4398_ _1106_ _0378_ _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_141_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8288__A3 _3385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7251_ _2381_ _2389_ _2390_ _2392_ _2393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_105_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6299__A2 _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6202_ _1453_ _1456_ _1459_ _1295_ _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_125_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7182_ _2331_ _2332_ _0161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7248__A1 _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6133_ _1372_ _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8445__B1 _3541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7799__A2 _2921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8996__A1 _3230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6064_ _1303_ _0886_ _1304_ _1305_ _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_112_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5015_ _4478_ _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7221__I as2650.addr_buff\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8748__A1 _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8599__I1 _3017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6223__A2 _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6966_ _2163_ _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8480__C _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7971__A2 _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7377__B _2403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8705_ _3792_ _3793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5917_ _0763_ _1105_ _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6897_ _2082_ _2088_ _2106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_70_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8636_ _3724_ _3725_ _3726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5848_ _0378_ _1071_ _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7723__A2 _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8920__A1 _3962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8567_ _0436_ _3481_ _3426_ _3652_ _3526_ _3661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_107_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5779_ _1039_ _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7518_ _2642_ _2647_ _2653_ _2502_ _2654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_135_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8498_ _0952_ _3561_ _3594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_108_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7449_ _1554_ _0358_ _2586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6300__I _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7239__A1 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9119_ _0012_ clknet_leaf_38_wb_clk_i as2650.stack\[5\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8987__A1 _3336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8227__I _3287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4755__I _4324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8739__A1 _3144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6214__A2 _4489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6970__I _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_48_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5973__A1 _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8911__A1 _3966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5725__A1 as2650.pc\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5725__B2 as2650.r123_2\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7478__A1 _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5535__B _4321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9240__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6150__A1 _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8565__C _3001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7650__A1 as2650.pc\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4665__I _4245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6453__A2 _1692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6820_ _2003_ _2011_ _2032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7953__A2 _2441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6751_ _1882_ _1965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5702_ as2650.pc\[11\] _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6682_ as2650.stack\[1\]\[8\] _1909_ _1910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5429__C _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8902__A1 _4153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8421_ as2650.stack\[0\]\[5\] _3361_ _3362_ as2650.stack\[1\]\[5\] _3520_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_5633_ as2650.pc\[4\] _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_117_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8352_ _3371_ _3452_ _3420_ _3453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5564_ _4215_ _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7303_ _4200_ _1364_ _1363_ _2442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_8283_ as2650.stack\[0\]\[2\] _3319_ _3320_ as2650.stack\[1\]\[2\] _3385_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_144_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5495_ as2650.holding_reg\[7\] _0799_ _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_144_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8130__A2 _3061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6120__I _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7234_ _1579_ _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6141__A1 _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8756__B _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6692__A2 _1909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7165_ _2175_ _2248_ _2322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8969__A1 _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6116_ _1377_ _4527_ _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7096_ _2269_ _0138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4575__I _4155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6444__A2 _1685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6047_ _4214_ _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8984__A4 _4023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8197__A2 _4180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9113__CLK clknet_leaf_67_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7998_ _3119_ _3120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_81_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6949_ _1500_ _1309_ _2154_ _2155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_35_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8619_ _1251_ _3709_ _3710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9263__CLK clknet_leaf_52_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6380__A1 _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8121__A2 _2155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6132__A1 _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7880__A1 _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6683__A2 _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6965__I _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6186__B _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4997__A2 _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7796__I _2925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6199__A1 _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5946__A1 _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6205__I _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7699__A1 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8360__A2 _3428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5174__A2 _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8112__A2 _3153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5280_ _0582_ _0584_ _0587_ _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__8663__A3 _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7871__A1 _2982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7871__B2 _2998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4685__A1 _4264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8970_ _1555_ _2634_ _4010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__9136__CLK clknet_leaf_58_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7921_ _3045_ _2354_ _3046_ _2433_ _3047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__4988__A2 _4332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8179__A2 _2435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7852_ net53 _2942_ _2943_ _2981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7926__A2 _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6803_ _1986_ _2015_ _2016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5937__A1 _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9286__CLK clknet_leaf_27_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7783_ _0964_ _0757_ _2913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4995_ _4290_ _4293_ _4302_ _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_71_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6734_ _0788_ _1736_ _1890_ _1948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_32_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6665_ _1886_ _1893_ _1894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_108_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5954__I _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8351__A2 _3425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7154__A3 _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8404_ _3221_ _3499_ _3502_ _1294_ _3503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_34_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5616_ _0917_ _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5165__A2 _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9384_ _0277_ clknet_leaf_3_wb_clk_i as2650.overflow vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6596_ _1800_ _1821_ _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_121_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8335_ _2793_ _3435_ _3076_ _3436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_121_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5547_ _0850_ _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8266_ _2391_ _3369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5478_ _0438_ _0782_ _0783_ _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__7862__A1 as2650.pc\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7217_ as2650.addr_buff\[2\] _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8197_ as2650.pc\[0\] _4180_ _3301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_132_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7148_ _1411_ _2307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7614__A1 net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8811__B1 _3847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7079_ _2258_ _2252_ _2253_ as2650.stack\[1\]\[2\] _2254_ _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_115_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8590__A2 _3665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout51 net25 net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7565__B _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8342__A2 _3425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5156__A2 _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6353__A1 _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6353__B2 _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7853__A1 _2521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9159__CLK clknet_leaf_58_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7605__A1 _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9070__A3 _4062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8030__A1 _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5919__A1 _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6187__A4 _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4780_ _4360_ _4361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5395__A2 _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5774__I _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8333__A2 _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6450_ _1502_ _1692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5147__A2 _4522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5401_ as2650.stack\[3\]\[13\] _4479_ _0427_ as2650.stack\[2\]\[13\] _0707_ _0708_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6381_ _4467_ _4463_ _1637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8120_ _3170_ _3230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5332_ _0638_ _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7844__A1 _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8051_ _3163_ _3164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5263_ _4502_ _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_130_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7844__B2 _2928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7002_ _2201_ _2164_ _2168_ as2650.stack\[2\]\[6\] _2173_ _2202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_69_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9046__B1 _4079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5194_ _0502_ _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8953_ _3995_ _2076_ _4000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7904_ _2963_ _3013_ _3030_ _3031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8325__I _2387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8884_ _3947_ _3949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4830__A1 _4354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7835_ _2960_ _2962_ _2963_ _2964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_110_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7766_ _2896_ _2897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5386__A2 _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4978_ _4348_ _0288_ _4506_ _4509_ _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_36_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5630__I0 _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6717_ _1672_ _1925_ _1932_ _0096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_20_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7697_ _1680_ _2588_ _2829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9436_ net46 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6648_ as2650.r0\[5\] _1745_ _1877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6335__A1 as2650.psu\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6335__B2 as2650.psu\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_9367_ _0260_ clknet_leaf_68_wb_clk_i as2650.r123\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6579_ _1809_ _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8088__A1 _2383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8318_ _3376_ _3420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9301__CLK clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9298_ _0191_ clknet_leaf_2_wb_clk_i as2650.holding_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8249_ _2335_ _3347_ _3351_ _3352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_106_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7404__I _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9037__B1 _3141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6464__B _1702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8563__A2 _3647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6169__A4 _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6574__A1 _4519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5621__I0 _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5594__I _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5129__A2 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6326__A1 _4463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6326__B2 _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6877__A2 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8838__C _3910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9015__B _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5301__A2 _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8251__A1 _1681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5950_ _1056_ _1223_ _1224_ _1053_ _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_94_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4812__A1 _4172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8003__A1 _3122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4901_ _4481_ _4482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5881_ as2650.r123_2\[0\]\[4\] _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_45_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7620_ _2154_ _2754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4832_ _4346_ _4353_ _4411_ _4412_ _4413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_107_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5368__A2 _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7551_ _1513_ _2686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_18_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4763_ _4343_ _4344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8306__A2 _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6502_ _0337_ _1736_ _1733_ _4441_ _1737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6317__A1 _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7482_ _2543_ _2603_ _2604_ _2619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4694_ _4274_ _4275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_53_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9221_ _0114_ clknet_leaf_37_wb_clk_i as2650.stack\[4\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6433_ _1674_ _1661_ _1675_ _0069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_106_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8748__C _3833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9152_ _0045_ clknet_leaf_16_wb_clk_i net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6364_ _1281_ _1615_ _1620_ _1611_ _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5540__A2 _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7817__A1 net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8103_ _3045_ _3214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5315_ as2650.stack\[3\]\[12\] _0622_ _4454_ _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6295_ _0373_ _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9083_ _4112_ _4115_ _3619_ _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_103_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7293__A2 _4237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8034_ _1626_ _3148_ _3149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5246_ _0544_ _0547_ _0552_ _0553_ _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_130_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5177_ _4269_ _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8793__A2 _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8936_ _3985_ _3986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8867_ _2294_ _3935_ _3938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7818_ _2945_ _2946_ _2947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_52_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6556__A1 _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8798_ _1627_ _0639_ _3880_ _3851_ _3881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_101_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7749_ _2876_ _2878_ _2880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7808__A1 _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8481__A1 _2645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5295__A1 _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5047__B2 _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8784__A2 _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6795__A1 _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5598__A2 _4466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9347__CLK clknet_leaf_40_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5538__B _4546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5770__A2 _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8568__C _3373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5100_ _0407_ _0310_ _0408_ _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_6080_ _1343_ _1352_ _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__8472__A1 _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7275__A2 _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7979__I _2793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5031_ _0341_ _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8224__A1 _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5720__C _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7027__A2 _4482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8224__B2 _3327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8775__A2 _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6982_ _0925_ _2176_ _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8721_ _3219_ _0422_ _3183_ _3806_ _3807_ _3808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5933_ _1206_ _1207_ _0555_ _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_50_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_80_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8527__A2 _3594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8652_ _2577_ _3742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5864_ _0533_ _1119_ _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_61_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7603_ _2736_ _4246_ _2737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4815_ _4154_ _4395_ _4396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8583_ _2481_ _2354_ _3676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5210__A1 _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5795_ _1064_ _1066_ _1075_ _1076_ _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_72_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6123__I _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7534_ _1594_ _2555_ _2662_ _2669_ _2670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4746_ _4322_ _4325_ _4326_ _4327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5761__A2 _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7465_ _2601_ _2602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4677_ as2650.ins_reg\[5\] _4158_ _4177_ _4258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_107_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9204_ _0097_ clknet_leaf_46_wb_clk_i as2650.stack\[0\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6416_ _1658_ _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6710__A1 as2650.stack\[0\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7396_ _1340_ _2533_ _2534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput17 net17 io_oeb[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput28 net28 io_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_89_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9135_ _0028_ clknet_leaf_58_wb_clk_i as2650.stack\[5\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput39 net39 io_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_6347_ net3 _1604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9066_ _4100_ _3128_ _3127_ _4101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6278_ _1535_ _0840_ _1536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8017_ _0579_ _2399_ _3135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5229_ _4439_ _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7018__A2 _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5029__A1 _4277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6226__B1 _1480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8919_ _0523_ _3959_ _3973_ _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_77_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_38_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8518__A2 _3596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7726__B1 _2688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5201__A1 _4533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6968__I _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6701__A1 _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5504__A2 _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7257__A2 _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5268__A1 _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_77_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8206__A1 _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5540__C _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6217__B1 _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8757__A2 _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5112__I _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5440__A1 _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4951__I _4530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7980__A3 _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5991__A2 _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7193__A1 _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4600_ _4180_ _4181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_5580_ as2650.cycle\[1\] _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5743__A2 _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5782__I _4377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7250_ _1486_ _2391_ _1702_ _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__8693__A1 _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6299__A3 _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6201_ _0824_ _1458_ _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7181_ _2307_ _2322_ _2332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7248__A2 _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8445__A1 _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6132_ _0579_ _1398_ _1400_ _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8445__B2 _3542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8996__A2 _4029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6063_ _1335_ _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5014_ as2650.stack\[4\]\[9\] _4481_ _4460_ as2650.stack\[6\]\[9\] _0324_ as2650.stack\[5\]\[9\]
+ _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_85_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8748__A2 _3780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7658__B _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6965_ _0912_ _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_41_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4861__I _4211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8704_ _2423_ _3792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_81_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7971__A3 _3095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5916_ as2650.r123_2\[0\]\[6\] _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_74_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6896_ _2073_ _2097_ _2098_ _2104_ _2105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_8635_ as2650.pc\[13\] _1002_ _0995_ _3663_ _3725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_74_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5847_ _1065_ _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8566_ _3658_ _3659_ _3660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5778_ _1041_ _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6931__A1 _1795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7517_ _2643_ _2532_ _2652_ _2653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4729_ _4256_ _4304_ _4308_ _4309_ _4310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_8497_ _0966_ _3374_ _3593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7448_ _0351_ _0357_ _0374_ _2585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_107_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5498__A1 _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7379_ _0865_ _2517_ _2465_ _2518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7239__A2 _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8436__A1 _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9118_ _0011_ clknet_leaf_39_wb_clk_i as2650.stack\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8987__A2 _4010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9049_ _0467_ _0476_ _4084_ _4085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_77_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7412__I _2549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6998__A1 _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9192__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8739__A2 _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6028__I _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5422__A1 _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5273__I1 as2650.r123\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5973__A2 _4423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7175__A1 _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8911__A2 _1738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6922__A1 _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5725__A2 _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6698__I _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__9074__I _4105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7478__A2 _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8675__A1 _4398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6150__A2 _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8978__A2 _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4946__I _4525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7650__A2 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6750_ _1961_ _1963_ _1964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_17_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5701_ _0963_ _0993_ _0994_ _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6681_ _1907_ _1909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7166__A1 _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8902__A2 _4491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8420_ as2650.stack\[3\]\[5\] _2215_ _3519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5632_ _0617_ _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5716__A2 _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8351_ _3426_ _3425_ _3444_ _3446_ _3451_ _3327_ _3452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_106_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5563_ _4214_ _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8102__B _3212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7302_ _2437_ _2438_ _2440_ _2441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8666__A1 _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8282_ as2650.stack\[2\]\[2\] _3322_ _3384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5494_ _4368_ _4371_ _4373_ _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_117_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8130__A3 _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7233_ _4357_ _2370_ _2376_ _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5017__I _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7164_ _2285_ _2318_ _2319_ as2650.stack\[0\]\[1\] _2320_ _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_101_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5461__B _4546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6115_ _1373_ _1385_ _1386_ _1302_ _0040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_119_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8969__A2 _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7095_ as2650.r123\[3\]\[0\] _2269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6046_ _1034_ _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8772__B _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5687__I _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7997_ _3116_ _3117_ _3118_ _3119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__4591__I _4163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6948_ _0895_ _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6879_ _2082_ _2088_ _2089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_35_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8618_ _3708_ _3705_ _3353_ _3709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8549_ _3620_ _3621_ _3643_ _3592_ _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__6380__A2 _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8409__A1 _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5340__B1 _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7880__A2 _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5643__A1 _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7396__A1 _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5597__I _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5946__A2 _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7699__A2 _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8896__A1 as2650.stack\[7\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6221__I _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8648__A1 _3214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7320__A1 _4398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7871__A2 _2504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4685__A2 _4265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9073__A1 _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4676__I _4256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5634__A1 as2650.stack\[5\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7920_ _1462_ _1327_ _3046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_67_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8179__A3 _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7851_ _0990_ _2522_ _2979_ _2940_ _2980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_63_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8584__B1 _3675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6802_ _1987_ _2014_ _2015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_58_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7782_ _2911_ _1586_ _2912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5937__A2 _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4994_ _0302_ _0304_ _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6733_ _1945_ _1946_ _1947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7139__A1 _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7139__B2 as2650.stack\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6664_ _1888_ _1892_ _1893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8403_ _2996_ _3496_ _3500_ _3501_ _3502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5615_ _0361_ _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_9383_ _0276_ clknet_leaf_3_wb_clk_i as2650.carry vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6595_ _1189_ _1714_ _1825_ _0081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7227__I _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8334_ _2494_ _3424_ _3433_ _2352_ _3434_ _3435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__8639__A1 _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5546_ _0849_ _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8767__B _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8265_ _3360_ _3364_ _3365_ _3367_ _3368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_5477_ _0752_ _0343_ _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7311__A1 _4442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7216_ _1104_ _2358_ _2364_ _0163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5322__B1 _4461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7862__A2 _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8196_ _1442_ _3297_ _3299_ _3300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5873__A1 _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7147_ _2305_ _2286_ _2287_ as2650.stack\[3\]\[7\] _2277_ _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__9064__A1 _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8811__A1 _2109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7078_ _0921_ _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6029_ _1226_ _1286_ _1300_ _1302_ _0038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xclkbuf_leaf_5_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_5_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_104_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5389__B1 _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5928__A2 _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_3_0_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout52 net40 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8878__A1 _2305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8878__B2 as2650.stack\[7\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9380__CLK clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7550__A1 _2190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6353__A2 _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6105__A2 _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5864__A1 _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9055__A1 _4072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7605__A2 _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8802__A1 _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8030__A2 _3144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5120__I _4469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xwrapped_as2650_90 io_oeb[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__6041__A1 _4235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8869__A1 _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5400_ _0706_ _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_70_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6380_ _1515_ _1633_ _1636_ _0055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_75_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_75_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7491__B _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5331_ _0582_ _0584_ _0587_ _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8050_ _0898_ _3163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7844__A2 _2513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5262_ _0569_ _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5855__A1 _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7001_ _0947_ _2201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__9046__A1 _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5193_ _0495_ _0497_ _0501_ _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__9046__B2 _4081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9253__CLK clknet_leaf_55_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8952_ _0524_ _3992_ _3993_ as2650.r123\[2\]\[3\] _3999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_55_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7903_ _2961_ _3015_ _3030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8883_ _3947_ _3948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4830__A2 _4361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7834_ _2895_ _2912_ _2963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_58_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7765_ _2890_ _2894_ _2607_ _2896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4977_ _4305_ _4306_ _0287_ _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__7780__A1 _2774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4594__A1 _4174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6716_ as2650.stack\[0\]\[13\] _1923_ _1932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7696_ _1617_ _0828_ _2827_ _2828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_32_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9435_ net47 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6647_ as2650.r0\[4\] _1762_ _1876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6335__A2 _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9366_ _0259_ clknet_leaf_68_wb_clk_i as2650.r123\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6578_ as2650.r123\[0\]\[5\] as2650.r123_2\[0\]\[5\] _4144_ _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8317_ _3329_ _3382_ _3419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8088__A2 _3192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5529_ _0833_ _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9297_ _0190_ clknet_leaf_3_wb_clk_i as2650.holding_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8248_ _3048_ _3348_ _3350_ _1696_ _3351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_105_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9037__A1 _1627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8179_ _4444_ _2435_ _3281_ _3282_ _3283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_87_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7599__A1 _2694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8260__A2 _1637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6271__A1 _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output31_I net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6023__A1 _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7771__A1 _2785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6326__A2 _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9126__CLK clknet_leaf_59_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7826__A2 _2952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6629__A3 _1858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9276__CLK clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9028__A1 _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8251__A2 _3353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4900_ _4464_ _4481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8003__A2 _3123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5880_ _1142_ _1055_ _1158_ _0033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_61_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4831_ _4262_ _4412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7762__A1 _2203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7550_ _2190_ _2655_ _2685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4762_ _4279_ _4311_ _4340_ _4342_ _4343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_109_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6501_ _1723_ _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7481_ _2542_ _2618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7514__A1 _2643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4693_ _4273_ _4274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9220_ _0113_ clknet_leaf_40_wb_clk_i as2650.stack\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6432_ as2650.stack\[2\]\[14\] _1659_ _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_128_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9151_ _0044_ clknet_leaf_15_wb_clk_i net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6363_ _1619_ _1281_ _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8102_ _3090_ _1231_ _3212_ _3213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5314_ _4452_ _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7817__A2 net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9082_ _4108_ _4114_ _4115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6294_ _4531_ _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5828__A1 _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8033_ _1710_ _1294_ _3148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9019__A1 _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5245_ _4336_ _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8490__A2 _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5176_ _0479_ _0484_ _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_29_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7240__I _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6253__A1 _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6284__C _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8935_ _4272_ _1612_ _3985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_71_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_28_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5896__S _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8866_ _0921_ _3931_ _3932_ as2650.stack\[7\]\[2\] _3933_ _3937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_38_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_5_0_wb_clk_i clknet_0_wb_clk_i clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_101_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7817_ net37 net36 _2885_ _2946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_24_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8797_ _0342_ _3557_ _3879_ _3880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8071__I _3183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9149__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7748_ _2866_ _2876_ _2878_ _2879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_61_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7505__A1 _2638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7679_ _1559_ _2560_ _2811_ _2565_ _2812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_123_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9299__CLK clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9349_ _0242_ clknet_leaf_51_wb_clk_i as2650.stack\[7\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7415__I _2469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8481__A2 _3574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7284__A3 _4425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_67_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6492__B2 _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6244__A1 _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5047__A2 _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8690__B _3778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7992__A1 _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5598__A3 _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4949__I _4528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4730__A1 _4303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8472__A2 _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8584__C _3676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5030_ _0339_ _0340_ _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_140_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8224__A2 _3317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7027__A3 _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6235__A1 _4550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6981_ _2183_ _2171_ _2172_ as2650.stack\[2\]\[3\] _2173_ _2184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_47_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7983__A1 _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5932_ _0796_ _0800_ _0798_ _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_65_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8720_ _3143_ _4527_ _3080_ _3807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8651_ _3292_ _3727_ _3740_ _3373_ _3741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5863_ as2650.r123_2\[0\]\[3\] _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_94_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7602_ _0684_ _2736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6404__I _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4814_ _4162_ _4393_ _4394_ _4395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_142_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8582_ _2368_ _2385_ _3441_ _3675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5794_ _1062_ _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5210__A2 _4545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7533_ _2469_ _2668_ _2669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4745_ _4303_ _4310_ as2650.psl\[3\] as2650.carry _4326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_72_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7464_ as2650.pc\[2\] net8 _2601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4676_ _4256_ _4257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9203_ _0096_ clknet_leaf_47_wb_clk_i as2650.stack\[0\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6415_ _0984_ _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7395_ _0896_ _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput18 net18 io_oeb[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_9134_ _0027_ clknet_leaf_56_wb_clk_i as2650.stack\[5\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput29 net29 io_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__4721__A1 _4296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6346_ _1578_ _1602_ _1603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9065_ _4072_ _4100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8463__A2 _3560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6277_ _4227_ _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8016_ _3120_ _3133_ _3134_ _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5228_ _4494_ _0534_ _0536_ _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_102_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5159_ _0393_ _0467_ _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_84_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5029__A2 _4423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6226__A1 _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6226__B2 _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7974__A1 net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8918_ _3962_ _1772_ _3964_ as2650.r123\[1\]\[3\] _3973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_71_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7726__A1 net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8849_ _3921_ _3922_ _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7726__B2 _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6314__I _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5201__A2 _4524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6701__A2 _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6984__I _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6217__A1 _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9314__CLK clknet_leaf_9_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6217__B2 _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6768__A2 _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4779__A1 _4333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8704__I _2423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5440__A2 _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6224__I _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7193__A2 _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8693__A2 _3766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6299__A4 _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6200_ _0754_ _1457_ _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7180_ _2305_ _2318_ _2319_ as2650.stack\[0\]\[7\] _2309_ _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_131_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6131_ _1399_ _0694_ _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7248__A3 _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8445__A2 _2777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5259__A2 _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6062_ net3 _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5013_ _4468_ _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_61_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5303__I _4348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6208__A1 _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7956__A1 _1617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6964_ _2138_ _2143_ _2169_ _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_81_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5431__A2 _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8703_ _0619_ _3368_ _3791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_74_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5915_ _1177_ _1160_ _1191_ _0035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_53_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6895_ _2093_ _2096_ _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8634_ as2650.pc\[14\] _3724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5846_ _1052_ _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_50_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8565_ _3250_ _3645_ _3651_ _2492_ _3001_ _3659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5777_ _1058_ _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_3_5_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7516_ _2648_ _2650_ _2651_ _1340_ _2652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_124_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4728_ _4291_ _4256_ _4309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_8496_ _0953_ _3289_ _3591_ _3592_ _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_33_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8133__A1 _3151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7447_ _2556_ _2582_ _2583_ _2584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_50_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4659_ _4238_ _4239_ _4165_ _4240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_107_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5498__A2 _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7378_ _1359_ _2517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6329_ _0755_ _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_9117_ _0010_ clknet_leaf_41_wb_clk_i as2650.stack\[5\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8436__A2 _2539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9337__CLK clknet_leaf_77_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9048_ _0561_ _0569_ _4082_ _4083_ _4084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_49_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7947__A1 _3069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5422__A2 _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8372__A1 _2648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6979__I _2181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5186__A1 _4521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6922__A2 _2129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4933__A1 _4511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8124__A1 _3230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8675__A2 _2632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6686__A1 _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5489__A2 _4376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5110__A1 _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8862__C _3933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7938__A1 _2824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_29_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_29_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_36_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4962__I _4541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5413__A2 _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5700_ as2650.stack\[6\]\[10\] _0986_ _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6680_ _1907_ _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8363__A1 _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5631_ _0931_ _0011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8350_ _3447_ _3448_ _3449_ _3450_ _3451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_5562_ _0850_ _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4924__A1 _4305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7301_ _4431_ _1256_ _2439_ _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_8281_ as2650.stack\[3\]\[2\] _4474_ _4473_ _3383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8666__A2 _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5493_ _0797_ _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_117_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7232_ _1706_ _2363_ _2376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8130__A4 _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7163_ _2309_ _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6429__A1 as2650.stack\[2\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6114_ net42 _1380_ _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7094_ _2267_ _2268_ _0137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_28_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6045_ _1314_ _1317_ _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5101__A1 _4277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6129__I _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7929__A1 _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5968__I _4427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7996_ _1277_ _1493_ _1517_ _0852_ _3118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_54_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6947_ _0881_ _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8354__A1 _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6878_ _2086_ _2087_ _2088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8617_ as2650.pc\[13\] _3707_ _3708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_139_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5829_ _1062_ _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4915__A1 as2650.r123\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8548_ _3292_ _3624_ _3642_ _3331_ _3643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_10_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8106__A1 _3211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8479_ _1599_ _1490_ _3575_ _3576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8409__A2 _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7093__A1 _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8290__B1 _3155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6840__A1 _2021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7579__B _2554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7396__A2 _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8593__A1 _3035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5099__B _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5159__A1 _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8896__A2 _3947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9018__C _3742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6659__A1 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7320__A2 _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9034__B _4070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9073__A2 _4106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5634__A2 _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7850_ _2958_ _2967_ _2973_ _2978_ _2979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_75_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8584__A1 _2495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8584__B2 _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6801_ _1989_ _2013_ _2014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_24_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5398__A1 as2650.stack\[6\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7781_ as2650.pc\[9\] _2911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_17_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4993_ as2650.holding_reg\[1\] _0301_ _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_63_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6732_ _1870_ _1895_ _1946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7936__C _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8336__A1 _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6663_ _1890_ _1891_ _1892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7508__I _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8402_ _0685_ _2539_ _2396_ _3501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6412__I _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5614_ _0916_ _0009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6594_ as2650.r123_2\[1\]\[5\] _1729_ _1824_ _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_9382_ _0275_ clknet_3_2_0_wb_clk_i as2650.psl\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8333_ _2368_ _1490_ _1508_ _2651_ _3434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5545_ _4448_ _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5028__I _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8264_ as2650.stack\[7\]\[1\] _3366_ _3322_ as2650.stack\[6\]\[1\] _4476_ _3367_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_105_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5476_ _4445_ _0781_ _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7311__A2 _2449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7215_ _2362_ _2363_ _2364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8195_ _2899_ _2755_ _1276_ _3298_ _3299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_7146_ _2204_ _2305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9064__A2 _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7077_ _2255_ _2257_ _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8811__A2 _3844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6028_ _1301_ _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8575__A1 _2950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5389__A1 _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7979_ _2793_ _3103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout53 net38 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8878__A2 _3931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6322__I _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7550__A2 _2655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7302__A2 _2438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5864__A2 _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9055__A2 _3113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8693__B _2629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8802__A2 _3856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_80 io_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_91 io_oeb[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6041__A2 _4241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8869__A2 _3931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7328__I _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6232__I _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5552__A1 _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5330_ as2650.holding_reg\[5\] _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5261_ _0396_ _0543_ _0564_ _0568_ _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__5304__A1 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7000_ _2199_ _2200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5192_ _0500_ _4141_ _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9046__A2 _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7998__I _3119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_44_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_110_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8951_ _3997_ _3998_ _0264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7902_ _2836_ _3026_ _3028_ _2720_ _2486_ _3029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA_clkbuf_leaf_18_wb_clk_i_I clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6280__A2 _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8882_ _3946_ _3947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8557__A1 _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7833_ _2961_ _2962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_36_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7764_ _2890_ _2894_ _2895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8309__A1 _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4976_ _4243_ _4347_ _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6715_ _1670_ _1925_ _1931_ _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_71_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5791__A1 _4398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7695_ _2798_ _2802_ _2826_ _2827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_71_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9434_ net47 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6646_ _0671_ _1731_ _1875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8580__I1 _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9365_ _0258_ clknet_3_4_0_wb_clk_i as2650.r123\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6577_ _1805_ _1806_ _1807_ _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_118_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8316_ _3336_ _3382_ _3390_ _3369_ _3417_ _3418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_117_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5528_ _4375_ _0832_ _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_105_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9296_ _0189_ clknet_leaf_11_wb_clk_i as2650.idx_ctrl\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6099__A2 _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7296__A1 _4233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8247_ _0911_ _1618_ _3349_ _3350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5459_ _0759_ _4532_ _0764_ _4231_ _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_79_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7835__A3 _2963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_57_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9037__A2 _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8178_ _1347_ _1363_ _3282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_82_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7129_ _2258_ _2286_ _2287_ as2650.stack\[3\]\[2\] _2288_ _2293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_75_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7599__A2 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8796__A1 _3844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8796__B2 _3847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6271__A2 _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8548__A1 _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7857__B _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output24_I net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7220__A1 _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7148__I _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7523__A2 _2606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8720__A1 _3143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6987__I _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7287__A1 _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7039__A1 _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8787__A1 _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8787__B2 _2630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8539__A1 _2526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5470__B1 _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7767__B _2751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4812__A3 _4175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7211__A1 _2334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4970__I _4232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4830_ _4354_ _4361_ _4410_ _4345_ _4411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_34_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5222__B1 _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4761_ _4341_ _4308_ _4279_ _4342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6500_ _1734_ _1735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8011__I0 _3129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7480_ _2609_ _2505_ _2508_ _1555_ _2616_ _2617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_14_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4692_ _4137_ _4272_ _4273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6431_ _1015_ _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9150_ _0043_ clknet_leaf_15_wb_clk_i net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6362_ _1618_ _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8101_ _3209_ _1507_ _3212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5313_ _0620_ _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__9220__CLK clknet_leaf_40_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6293_ _1550_ _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_9081_ _4113_ _4100_ _3133_ _4114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7817__A3 _2885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5306__I _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5244_ _0548_ _0504_ _0551_ _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8032_ _3147_ _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9019__A2 _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5175_ _0348_ _0482_ _0483_ _0353_ _0370_ _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_60_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8778__A1 _3810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9370__CLK clknet_leaf_76_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7450__A1 _2585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6253__A2 _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8934_ _0846_ _3959_ _3984_ _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8865_ _3934_ _3936_ _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_77_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5976__I _4417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7202__A1 _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4880__I _4460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7816_ net53 _2945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_51_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8796_ _3844_ _2084_ _3878_ _3847_ _3777_ _3879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__8950__A1 _3995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7747_ _2703_ _2877_ _2878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_75_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5764__A1 _4223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4959_ _4515_ _4527_ _4537_ _4538_ _4539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_71_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7678_ _2473_ _2810_ _2811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5516__A1 _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6629_ _1827_ _1833_ _1858_ _1859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_137_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9348_ _0241_ clknet_leaf_41_wb_clk_i as2650.stack\[7\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7269__A1 _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9279_ _0172_ clknet_3_3_0_wb_clk_i net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5216__I _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6492__A2 _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8769__A1 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7441__A1 _2521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6244__A2 _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6047__I _4214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8690__C _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7992__A2 _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7744__A2 _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8941__A1 _3966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5755__A1 _4143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5507__A1 _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8211__B _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9243__CLK clknet_leaf_55_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8457__B1 _1656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4730__A2 _4310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9042__B _4070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7341__I _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6235__A2 _4341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6980_ _2182_ _2183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5931_ _0724_ _0797_ _0794_ _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8650_ _3738_ _3739_ _3526_ _3740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5862_ _1123_ _1055_ _1141_ _0032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_62_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8932__A1 _3976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7601_ _1180_ _0668_ _2734_ _2735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__5746__A1 as2650.stack\[5\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4813_ _4186_ _4394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8581_ _3533_ _3673_ _3674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5793_ _0301_ _1068_ _1069_ _1074_ _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_124_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7532_ _2665_ _2667_ _2668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4744_ _4192_ _4324_ _4325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7463_ _2591_ _2599_ _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4675_ _4181_ _4255_ _4256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__8121__B _3221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9202_ _0095_ clknet_leaf_47_wb_clk_i as2650.stack\[0\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6414_ _1653_ _1660_ _1662_ _0063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7394_ _2531_ _2532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput19 net19 io_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_9133_ _0026_ clknet_leaf_53_wb_clk_i as2650.stack\[5\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4721__A2 _4299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6345_ _1597_ _1598_ _1600_ _1601_ _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_116_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8999__A1 _3189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9064_ _1518_ _0801_ _4099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6276_ _1523_ _1524_ _1529_ _1533_ _1534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_115_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5227_ _0535_ _0343_ _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8015_ _0461_ _3120_ _3134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5158_ _0466_ _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7423__A1 _4390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6226__A2 _4187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5089_ as2650.holding_reg\[2\] _0355_ _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_44_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7974__A2 _3090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8917_ _3971_ _3972_ _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5985__A1 _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8082__I _1685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8848_ _2307_ _3912_ _3922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7726__A2 _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8923__A1 _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_77_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8779_ as2650.psl\[5\] _3792_ _3863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9266__CLK clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5201__A3 _4510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8687__B1 _4435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4960__A2 _4514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6330__I _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6162__A1 _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6701__A3 _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7161__I _2312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7414__A1 _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6217__A2 _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7414__B2 _2550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4779__A2 _4359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7193__A3 _4253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6528__I0 as2650.r123\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6240__I _1497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6130_ _1375_ _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4695__I _4262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6061_ _1318_ _1333_ _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7653__A1 _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7071__I _2246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9139__CLK clknet_leaf_46_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5012_ _0286_ _0293_ _0322_ _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7405__A1 as2650.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8602__B1 _3693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7939__C _2578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7956__A2 _2352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5967__A1 _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6963_ _2147_ _2164_ _2168_ as2650.stack\[2\]\[0\] _2142_ _2169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__8116__B _3220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6415__I _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8702_ _4227_ _3790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5914_ _1124_ _1179_ _1190_ _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__5459__C _4231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6894_ _2090_ _2092_ _2103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8905__A1 _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8633_ _3703_ _3723_ _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5845_ _0436_ _1088_ _1090_ _0437_ _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_139_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8564_ _3458_ _3645_ _3657_ _3391_ _3658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5776_ _1039_ _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7515_ _0508_ _1489_ _2651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4727_ _4305_ _4306_ _4307_ _4308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_8495_ _2577_ _3592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7246__I _2387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8133__A2 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7446_ _2581_ _0289_ _0291_ _2583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_68_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4658_ as2650.cycle\[5\] as2650.cycle\[4\] _4239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_107_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7892__A1 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6695__A2 _1907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7377_ _2490_ _2515_ _2403_ _2516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4589_ _4167_ _4169_ _4170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9116_ _0009_ clknet_leaf_42_wb_clk_i as2650.stack\[5\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6328_ _1584_ _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9047_ _0421_ _0451_ _0467_ _0475_ _4083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_49_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6259_ _1516_ _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7947__A2 _3071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5958__A1 _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6325__I _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5273__I3 as2650.r123_2\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8372__A2 _3469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5186__A2 _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7580__B1 _2709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4933__A2 _4512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8124__A2 _3231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7883__A1 _2982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6686__A2 _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4697__A1 _4159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7635__A1 _2752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5404__I _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5110__A2 _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7938__A2 _3063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8060__A1 _3154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5949__A1 _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_69_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_69_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7775__B _2550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8363__A2 _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5630_ _0925_ _0930_ _0860_ _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_32_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5561_ _0864_ _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4924__A2 _4306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7300_ _4423_ _1257_ _2439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_144_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8280_ _3381_ _3382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5492_ _0737_ _0732_ _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7874__A1 _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7231_ _4355_ _2370_ _2375_ _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7874__B2 _3001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4688__A1 _4233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7162_ _2315_ _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7626__A1 _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6429__A2 _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6113_ _1382_ _1376_ _1384_ _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7093_ _0951_ _2256_ _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5314__I _4452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6044_ _1316_ _1267_ _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_112_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5101__A2 _4324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7929__A2 _2453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7995_ _1457_ _1477_ _1571_ _3117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6145__I _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6946_ _1335_ _2151_ _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_35_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6877_ _4367_ _1812_ _2087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8354__A2 _3289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8616_ _3035_ _3687_ _3707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5828_ _0400_ _1103_ _1066_ _1108_ _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5168__A2 _4505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8547_ _3640_ _3641_ _3329_ _3642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5759_ _4157_ _4242_ _4245_ _1040_ _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_136_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6117__A1 _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8478_ _2153_ _1489_ _3575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9304__CLK clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6668__A2 _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5933__B _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7429_ _2559_ _2566_ _2567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4679__A1 _4254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8290__A1 _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7093__A2 _2256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8290__B2 _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4851__A1 _4312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8042__A1 _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4603__A1 _4155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5651__I0 _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8270__I _3287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5159__A2 _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6356__A1 _1611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8203__C _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7856__A1 _2982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6659__A2 _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7320__A3 _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9058__B1 _4093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7608__A1 _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5095__A1 _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8033__A1 _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8584__A2 _3665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6800_ _1996_ _1999_ _2012_ _2013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_24_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7780_ _2774_ _2909_ _2910_ _0181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5398__A2 _4461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6595__A1 _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7792__B1 _2921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4992_ _0302_ _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6731_ _1873_ _1894_ _1945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8336__A2 _3425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6662_ _4366_ _1720_ _1891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7544__B1 _2633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9327__CLK clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8401_ _4265_ _3157_ _3500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5613_ _0908_ _0914_ _0915_ _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_9381_ _0274_ clknet_leaf_44_wb_clk_i as2650.psu\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6593_ _1795_ _1823_ _1824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5309__I _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8332_ _1708_ _2641_ _3432_ _3433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5544_ _4295_ _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7952__C _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8263_ _1918_ _3366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5475_ _0776_ _0777_ _0780_ _0526_ _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_69_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7214_ _2357_ _2363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8194_ _4392_ _2410_ _3298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5322__A2 _4479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_47_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7145_ _2200_ _2279_ _2304_ _0152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8272__A1 _3333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7076_ _0908_ _2256_ _2257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_87_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6027_ _4438_ _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8024__A1 _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8575__A2 _3610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5389__A2 _4547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7978_ _3087_ _3101_ _3102_ _2578_ _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6929_ _2131_ _2132_ _2135_ _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_126_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout54 net35 net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7838__A1 _2923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7302__A3 _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7066__A2 _1905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5077__A1 _4359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8015__A1 _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_70 io_oeb[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_81 io_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_45_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_as2650_92 io_oeb[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_2673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5001__A1 _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5552__A2 _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7829__A1 _2613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5260_ _0565_ _0567_ _0396_ _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5191_ _0499_ _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8254__A1 _3355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5068__A1 _4525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8950_ _3995_ _2048_ _3998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4815__A1 _4154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7901_ net52 _3027_ _3028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_3_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8881_ _1019_ _3899_ _3946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8557__A2 _2976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7832_ as2650.pc\[9\] _0964_ _0756_ _2961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_64_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6568__A1 _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7763_ _2729_ _2727_ _2891_ _2893_ _2894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_4975_ _4501_ _4513_ _4549_ _0285_ _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__8309__A2 _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6714_ as2650.stack\[0\]\[12\] _1927_ _1931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5467__C _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7694_ _2825_ _0749_ _2826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9433_ net46 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6645_ _1844_ _1848_ _1874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9364_ _0257_ clknet_leaf_73_wb_clk_i as2650.r123\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6576_ _0363_ _1748_ _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8315_ _3391_ _3398_ _3414_ _2345_ _3416_ _3417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_117_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_3_wb_clk_i_I clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5527_ _0760_ _0761_ _0717_ _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_9295_ _0188_ clknet_leaf_11_wb_clk_i as2650.idx_ctrl\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7254__I _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6099__A3 _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8246_ _1679_ _2545_ _3349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8493__A1 _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5458_ _0598_ _0763_ _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8177_ _1322_ _0889_ _3279_ _3280_ _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_99_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5389_ _0670_ _4547_ _0693_ _0695_ _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_8_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8245__A1 _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7128_ _2289_ _2292_ _0147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5059__A1 _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8796__A2 _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7059_ as2650.r123_2\[3\]\[7\] _2242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8548__A2 _3624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7220__A2 _2358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output17_I net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8720__A2 _4527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5534__A2 _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8484__A1 _3415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7287__A2 _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5298__A1 _4378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5613__S _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8236__A1 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8787__A2 _2633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9172__CLK clknet_leaf_60_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6952__B _2155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8539__A2 _3623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5470__B2 as2650.stack\[6\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8723__I _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7211__A2 _2358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4760_ _4183_ _4225_ _4341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8011__I1 _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4691_ _4154_ _4189_ _4271_ _4272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8711__A2 _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6430_ _1672_ _1661_ _1673_ _0068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_70_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6361_ _1617_ _1618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8100_ _2386_ _3090_ _1370_ _3211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5312_ _0619_ _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8475__A1 _2925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9080_ _1622_ _4113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7007__C _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6292_ _1549_ _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8031_ _3146_ _0730_ _3130_ _3147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5243_ _0549_ _0550_ _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9019__A3 _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5174_ _4524_ _0290_ _0462_ _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_111_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8778__A2 _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8933_ as2650.r123\[1\]\[7\] _3964_ _3983_ _3984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_83_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5461__A1 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8864_ _2290_ _3935_ _3936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7815_ _2774_ _2941_ _2944_ _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7202__A2 _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8795_ net27 _1525_ _3792_ _3878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7249__I _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5213__A1 _4345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6153__I _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7746_ _1604_ _0829_ _2877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_40_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4958_ _4221_ _4538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5764__A2 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8789__B _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7677_ _2806_ _2809_ _2810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4889_ _4469_ _4470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6628_ _1836_ _1857_ _1858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_137_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6713__A1 _1668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5516__A2 _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7910__B1 _2507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9347_ _0240_ clknet_leaf_40_wb_clk_i as2650.stack\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6559_ _1774_ _1775_ _1790_ _1791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__7269__A2 _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9278_ _0171_ clknet_leaf_20_wb_clk_i net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5941__B _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8229_ _0865_ _3289_ _3332_ _3112_ _0208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9195__CLK clknet_leaf_47_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8769__A2 _2633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6328__I _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5232__I as2650.r123\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7587__C _2721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5388__B _4546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5204__A1 _4396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6063__I _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8941__A2 _1979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6952__A1 _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5755__A2 _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8699__B _3080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6180__A2 _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8457__A1 as2650.stack\[4\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8457__B2 as2650.stack\[5\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7622__I _2755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8209__A1 _3293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6235__A3 _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5930_ as2650.r123_2\[0\]\[7\] _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_47_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5861_ _1124_ _1125_ _1140_ _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__7196__A1 _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7600_ _2663_ _2732_ _2710_ _2733_ _2734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__8932__A2 _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4812_ _4172_ _4166_ _4175_ _4393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_8580_ _0996_ _3006_ _0837_ _3673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_72_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5746__A2 _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5792_ _4392_ _1071_ _1073_ _1067_ _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_72_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7531_ _2584_ _2585_ _2666_ _2667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4743_ _4323_ _4178_ _4324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8402__B _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7462_ _1555_ _2560_ _2597_ _2598_ _2599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__8696__A1 _3703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4674_ as2650.ins_reg\[3\] _4255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_9201_ _0094_ clknet_leaf_60_wb_clk_i as2650.stack\[0\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6413_ as2650.stack\[2\]\[8\] _1661_ _1662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7393_ _2153_ _2384_ _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_134_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9132_ _0025_ clknet_leaf_56_wb_clk_i as2650.stack\[5\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8448__A1 _3459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6344_ _1238_ _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_1_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4721__A3 _4301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_9063_ _1212_ _1431_ _4098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6275_ _1273_ _1456_ _1531_ _1532_ _1533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_88_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8014_ _0535_ _1295_ _3132_ _3133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5226_ _0492_ _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5052__I as2650.r0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5157_ _0461_ _0314_ _0465_ _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8620__A1 _2996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5987__I _4369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5088_ as2650.holding_reg\[2\] _0355_ _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_42_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7974__A3 _2155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8916_ _0424_ _3969_ _3972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7187__A1 _2336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8847_ _2305_ _3908_ _3909_ as2650.stack\[6\]\[7\] _3900_ _3921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8384__B1 _1656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5001__B _4325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8923__A2 _1939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8778_ _3810_ _0694_ _3862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7729_ _2850_ _2853_ _2860_ _1450_ _2861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_40_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6611__I _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8687__A1 _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8439__A1 _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9100__A2 _4129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7111__A1 _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7442__I _2520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8611__A1 _3035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7178__A1 _2265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9210__CLK clknet_leaf_77_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5728__A2 _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7617__I _2483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_15_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9360__CLK clknet_leaf_59_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6528__I1 as2650.r123_2\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7350__A1 _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8876__C _3933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7653__A2 _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6060_ _1319_ _1321_ _1332_ _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_112_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input8_I io_in[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5011_ _0296_ _0321_ _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7405__A2 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8602__A1 _3082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8602__B2 _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7301__B _2439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6962_ _2167_ _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5600__I _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5913_ _1126_ _1189_ _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8701_ _1552_ _1541_ _3170_ _3789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6893_ _1174_ _1938_ _2102_ _0102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7169__A1 _2294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8632_ _1008_ _3377_ _3722_ _3723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5844_ _1053_ _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6916__A1 _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8563_ _3504_ _3647_ _3649_ _3459_ _3103_ _3656_ _3657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_33_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5775_ _1041_ _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7514_ _2643_ _2649_ _2650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4726_ as2650.holding_reg\[0\] _4307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8494_ _3333_ _3563_ _3590_ _3591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7445_ _0289_ _0291_ _2581_ _2582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6144__A2 _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4657_ as2650.cycle\[6\] _4238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7892__A2 _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7376_ _2145_ _2496_ _2512_ _2513_ _2514_ _2515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_4588_ as2650.cycle\[1\] _4168_ _4169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9115_ _0008_ clknet_leaf_38_wb_clk_i as2650.stack\[5\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6327_ net9 _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8358__I _3393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9094__A1 _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9046_ _0421_ _0451_ _4079_ _4081_ _4082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_67_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8841__A1 _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6258_ _1095_ _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5209_ _0517_ _4526_ _4545_ _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_76_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6189_ _4311_ _1445_ _1446_ _1447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_44_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5407__A1 _4274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9233__CLK clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7211__B _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5958__A2 _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9383__CLK clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7580__A1 _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7580__B2 _4268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5385__C _4378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6135__A2 _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7332__A1 _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7883__A2 _2942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5894__A1 _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8268__I _3290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9085__A1 _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8832__A1 _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5621__S _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7399__A1 _2530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4745__B as2650.psl\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5949__A2 _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6071__A1 _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8899__A1 _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7020__B1 _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7347__I _2485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7571__A1 _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6251__I _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5560_ _0863_ _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4924__A3 _4503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_38_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_89_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5491_ _0721_ _0723_ _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7230_ _1292_ _2359_ _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4700__S _4147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7874__A2 _2525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4688__A2 _4206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_37_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7161_ _2312_ _2318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__9076__A1 _3138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6112_ _1377_ _1383_ _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7626__A2 _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7092_ _2205_ _2252_ _2253_ as2650.stack\[1\]\[7\] _2243_ _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_86_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5637__A1 _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9256__CLK clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6043_ _1315_ _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_98_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7810__I _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7994_ _1367_ _2420_ _3116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6945_ _2150_ _4176_ _2151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8641__I _3081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9000__A1 _3492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6876_ _2083_ _2085_ _2086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_35_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8615_ _3705_ _3706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5827_ _1104_ _1105_ _1107_ _1068_ _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7562__A1 _2636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_76_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8546_ _0335_ _3369_ _3317_ _3624_ _3641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5758_ _4149_ _4198_ _4151_ _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__8797__B _3879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4709_ _4190_ _4283_ _4289_ _4290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_8477_ _1679_ _2849_ _3573_ _3574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7314__A1 _2406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5689_ _0979_ _0980_ _0973_ as2650.r123_2\[0\]\[1\] _0983_ _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_108_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7428_ _2536_ _2560_ _2563_ _2565_ _2566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5876__A1 _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4679__A2 _4259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7206__B _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7359_ _2418_ _1710_ _2497_ _2498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9067__B2 _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8814__A1 _2630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5628__A1 as2650.stack\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9029_ _4365_ _1251_ _4066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4851__A2 _4431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8042__A2 _2461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6053__A1 _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4603__A2 _4183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5651__I1 as2650.stack\[5\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6356__A2 _1612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9129__CLK clknet_leaf_58_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7305__A1 _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5867__A1 _4188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9279__CLK clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9058__A1 _4089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9058__B2 _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5331__A3 _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5415__I _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7608__A2 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8281__A2 _4474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5095__A2 _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4842__A2 _4278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8033__A2 _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6044__A1 _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4991_ as2650.holding_reg\[1\] _0301_ _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7792__A1 _2836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7792__B2 _2720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6730_ _1865_ _1897_ _1943_ _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6661_ _1807_ _1876_ _1889_ _1846_ _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__7544__A1 _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8400_ _0939_ _1614_ _3498_ _3499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5612_ _0859_ _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_9380_ _0273_ clknet_leaf_44_wb_clk_i as2650.psu\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6592_ _1798_ _1822_ _1823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_118_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8331_ _2182_ _1617_ _3432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5543_ _0786_ _4440_ _0793_ _0847_ _0007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8262_ as2650.stack\[4\]\[1\] _3361_ _3362_ as2650.stack\[5\]\[1\] _3365_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_144_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5474_ as2650.stack\[3\]\[14\] _4478_ _0527_ as2650.stack\[2\]\[14\] _0779_ _0780_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_121_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5858__A1 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7213_ _2361_ _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9049__A1 _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8193_ _1695_ _3295_ _3296_ _1509_ _3297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_113_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7144_ _2265_ _2281_ _2283_ as2650.stack\[3\]\[6\] _2288_ _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_119_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8272__A2 _3335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7075_ _2175_ _2166_ _2256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7480__B1 _2508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6026_ _1287_ _1299_ _1286_ _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_39_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4833__A2 _4344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8024__A2 _3140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6035__A1 _4263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7977_ net51 _3087_ _3102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5995__I _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5928__C _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6928_ _2133_ _2134_ _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7535__A1 _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6859_ _2058_ _2069_ _2070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_35_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8529_ _3623_ _3624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5849__A1 _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8974__C _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5077__A2 _4525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8015__A2 _3120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6026__A1 _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_60 io_oeb[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_3386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7774__A1 _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_as2650_71 io_oeb[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xwrapped_as2650_82 io_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__4588__A1 as2650.cycle\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_as2650_93 io_oeb[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4760__A1 _4183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5190_ _0498_ _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4815__A2 _4395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7900_ net39 _2983_ _3027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8880_ _3944_ _3945_ _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_64_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7831_ _2959_ _2960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6704__I _1923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7762_ _2203_ _0755_ _2892_ _2893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4974_ _0284_ _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_53_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_53_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6713_ _1668_ _1924_ _1930_ _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_71_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7517__A1 _2643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7693_ _0756_ _2825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_127_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9432_ net46 net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6644_ _1871_ _1855_ _1872_ _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6575_ _0498_ _1731_ _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9363_ _0256_ clknet_leaf_69_wb_clk_i as2650.r123\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_30_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8314_ _3415_ _3382_ _3409_ _2549_ _2856_ _3416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5526_ _4408_ _0830_ _0700_ _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_9294_ _0187_ clknet_leaf_25_wb_clk_i net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8245_ _1696_ _3334_ _1276_ _3348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_105_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5457_ _0679_ _0762_ _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6099__A4 _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8176_ _2156_ _2506_ _1364_ _4200_ _3280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5388_ _0517_ _0694_ _4546_ _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7127_ _2290_ _2291_ _2292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7270__I _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6256__A1 _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5059__A2 _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7058_ _2241_ _0128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6009_ _1282_ _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_74_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6008__A1 _4214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7756__A1 _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4990__A1 _4381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8181__A1 _3157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5298__A2 _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8236__A2 _4281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6247__A1 _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9317__CLK clknet_leaf_25_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7995__A1 _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6952__C _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7747__A1 _2703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8795__I0 net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5222__A2 _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4981__A1 _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4690_ _4213_ _4222_ _4231_ _4270_ _4271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_53_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8172__A1 _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4979__I _4508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7355__I _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6722__A2 _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6360_ _1616_ _1617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5311_ _0618_ _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6291_ _4391_ _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8475__A2 _3163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8030_ _1530_ _3144_ _3145_ _3146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_130_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5242_ _4332_ _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8186__I _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5173_ _4509_ _0481_ _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_60_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6238__A1 _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8119__C _3229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7986__A1 _3107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6789__A2 _2001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput1 io_in[10] net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_84_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8932_ _3976_ _1898_ _3983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_42_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5461__A2 _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8863_ _0968_ _2314_ _3935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6434__I _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7814_ _2919_ _2942_ _2943_ _2944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8794_ _3838_ _0740_ _3184_ _3875_ _3876_ _3877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_101_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5213__A2 _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7745_ _2806_ _2809_ _2875_ _2831_ _2876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_61_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4957_ _4531_ _4532_ _4536_ _4231_ _4537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_33_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4972__A1 _4551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7676_ _2807_ _2741_ _2808_ _2809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_4888_ _4468_ _4469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8163__A1 _4176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4889__I _4469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6627_ _1837_ _1856_ _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7910__A1 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7910__B2 _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6558_ _1779_ _1787_ _1789_ _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_9346_ _0239_ clknet_leaf_37_wb_clk_i as2650.stack\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5509_ _0447_ _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9277_ _0170_ clknet_leaf_20_wb_clk_i net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6489_ _0294_ _4152_ _4419_ _1236_ _1725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_8228_ _0865_ _3292_ _3330_ _3331_ _3332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_105_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8096__I _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8159_ _3263_ _3074_ _1511_ _3264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_59_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5513__I _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6229__A1 _4551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7977__A1 net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7729__B2 _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6344__I _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6401__A1 _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5204__A2 _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6952__A2 _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8154__A1 _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7901__A1 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4715__A1 _4295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8457__A2 _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5851__C _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5860_ _1126_ _1139_ _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7196__A2 _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8393__A1 _3492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7794__B _2922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4811_ _4391_ _4392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_61_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5791_ _4398_ _1072_ _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7530_ _0374_ _0351_ _0357_ _2666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_4742_ _4160_ _4323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7461_ _2564_ _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4673_ _4163_ _4253_ _4254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9200_ _0093_ clknet_leaf_60_wb_clk_i as2650.stack\[0\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6412_ _1659_ _1661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7392_ net29 _2530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9131_ _0024_ clknet_leaf_49_wb_clk_i as2650.stack\[5\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6343_ as2650.psl\[7\] _1599_ _1581_ _4248_ _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__8909__I _3961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7813__I _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9062_ _4064_ _4095_ _4096_ _4097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6274_ _4418_ _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5225_ _4485_ _0533_ _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8013_ _1594_ _1622_ _3132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7969__B _2508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5156_ _0314_ _0464_ _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7959__A1 _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4890__B1 _4470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8081__B1 _3067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8620__A2 _3705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5087_ _4341_ _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_56_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8915_ _3966_ _1753_ _3967_ as2650.r123\[1\]\[2\] _3971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_37_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8580__S _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8846_ _2199_ _3902_ _3920_ _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7187__A2 _4241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8777_ _3838_ _0662_ _3184_ _3859_ _3860_ _3861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__6934__A2 _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5989_ _0874_ _4330_ _1262_ _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7728_ _2204_ _2496_ _2859_ _2860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7659_ _1619_ _2790_ _2791_ _2792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8687__A2 _3769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9162__CLK clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8439__A2 _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9329_ _0222_ clknet_3_6_0_wb_clk_i as2650.pc\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7111__A2 _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8611__A2 _3374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5425__A2 _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8375__A1 _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_56_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8127__A1 _3081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7350__A2 _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_27_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_4_0_wb_clk_i clknet_0_wb_clk_i clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_113_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5010_ _0320_ _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8602__A2 _3686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6613__A1 _4382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5416__A2 _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6961_ _2165_ _2166_ _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5967__A3 _4432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5102__B _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8700_ _3219_ _0321_ _3183_ _3786_ _3787_ _3788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_81_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5912_ _0662_ _1188_ _1082_ _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__8366__A1 _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6892_ as2650.r123_2\[2\]\[4\] _1942_ _2101_ _2102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_74_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8631_ _3379_ _3720_ _3721_ _3420_ _3722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__8905__A3 _3958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5843_ as2650.r123_2\[0\]\[2\] _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6916__A2 _2109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5719__A3 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8562_ _3533_ _3651_ _3655_ _3656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_66_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9185__CLK clknet_leaf_73_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5774_ _1052_ _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7513_ net30 net29 net28 _2649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4725_ _4289_ _4306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8493_ _3371_ _3589_ _3376_ _3590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5328__I as2650.r123\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7444_ net7 _2581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4656_ _4236_ _4237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5352__A1 _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7375_ _1374_ _2514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4587_ as2650.cycle\[0\] _4168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_115_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9114_ _0007_ clknet_leaf_67_wb_clk_i as2650.r123\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6326_ _4463_ _1104_ _0375_ _0849_ _1583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_116_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9094__A2 _4113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9045_ _4335_ _4080_ _4081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6257_ _1475_ _1485_ _1512_ _1514_ _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__5063__I net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5208_ _4212_ _0516_ _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_76_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6188_ _1252_ _0403_ _0720_ _0801_ _1446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_69_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5998__I _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5139_ _0447_ _4314_ _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5407__A2 _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6604__A1 _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_8_wb_clk_i clknet_3_3_0_wb_clk_i clknet_leaf_8_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_44_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6080__A2 _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8829_ _3905_ _3909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8109__A1 _3219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5591__A1 _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5343__A1 _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6540__B1 _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5894__A2 _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9085__A2 _4113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8832__A2 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8284__I _1637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9320__D _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7399__A2 _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8596__A1 _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4745__C as2650.carry vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8217__C _4475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8060__A3 _3165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6071__A2 _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8348__B2 as2650.stack\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4761__B _4279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8899__A2 _3949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7020__A1 _2147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7020__B2 as2650.stack\[4\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7571__A2 _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5490_ _0794_ _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_8_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8520__A1 _3426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7323__A2 _2438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5185__I1 as2650.r123\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4688__A3 _4268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7160_ _0848_ _2311_ _2317_ _0154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_125_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7087__A1 _2197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6111_ _4387_ _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7087__B2 as2650.stack\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7091_ _2200_ _2245_ _2266_ _0136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6042_ _4232_ _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7312__B _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6707__I _1922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8587__A1 _3153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7993_ _3113_ _3114_ _3115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6944_ _0868_ _2150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_54_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8339__A1 _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__9000__A2 _3122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6875_ _0750_ _2084_ _2085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6442__I _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8614_ as2650.pc\[13\] _3704_ _3705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_126_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5826_ _1106_ _1071_ _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5022__B1 _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8545_ _3637_ _3639_ _3640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5757_ _4407_ _1037_ _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4708_ _4288_ _4289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8476_ _0953_ _1605_ _3573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5688_ _4497_ _0981_ _0982_ _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7314__A2 _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4897__I _4450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7427_ _2564_ _2565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5325__A1 _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5325__B2 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4639_ _4214_ _4219_ _4220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_135_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5876__A2 _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7358_ _1545_ _2487_ _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5007__B _4338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9200__CLK clknet_leaf_60_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6309_ _1525_ _1515_ _1566_ _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8814__A2 _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7289_ _1230_ _2427_ _1350_ _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9028_ _0855_ _4017_ _4065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_76_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8578__A1 _3392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7250__A1 _1486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6053__A2 _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7002__A1 _2201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6356__A3 _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8750__A1 _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7892__B _2852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7305__A2 _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9315__D _0208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4600__I _4180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5867__A2 _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7069__A1 _2147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7069__B2 as2650.stack\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7608__A3 _2741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8805__A2 _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6816__A1 _2027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8569__A1 _2969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6044__A2 _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4990_ _4381_ _4385_ _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7792__A2 _2918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6262__I _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6660_ _0498_ _1748_ _1783_ _0362_ _1889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7544__A2 _2630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5611_ _0912_ as2650.stack\[5\]\[1\] _0913_ _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6591_ _1800_ _1821_ _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_121_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8330_ _3428_ _3429_ _3430_ _3431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5542_ _4275_ _0846_ _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_34_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8189__I _3095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6504__B1 _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5473_ _0778_ _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8261_ as2650.stack\[0\]\[1\] _3361_ _3362_ as2650.stack\[1\]\[1\] _3363_ _3364_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__9223__CLK clknet_leaf_40_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6211__B _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7212_ as2650.addr_buff\[1\] _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8192_ _2144_ _1695_ _3296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9049__A2 _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7143_ _2193_ _2279_ _2303_ _0151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_98_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9373__CLK clknet_leaf_74_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7074_ _2170_ _2252_ _2253_ as2650.stack\[1\]\[1\] _2254_ _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_63_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7480__A1 _2609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6437__I _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6025_ _1290_ _1298_ _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7480__B2 _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7232__A1 _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8652__I _2577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7976_ _1692_ _3100_ _2403_ _3101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7783__A2 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8980__A1 _2342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5497__B _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6927_ _0752_ _2084_ _2126_ _2134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7268__I _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6858_ _2066_ _2068_ _2069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__7535__A2 _2592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8732__A1 _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5809_ _4295_ _0621_ _1085_ _1088_ _1090_ _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_126_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8601__B _3470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6789_ _1962_ _2001_ _2002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_13_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8528_ _3620_ _3622_ _3623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8099__I _3046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8459_ _3556_ _3557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8248__B1 _3350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8799__A1 _3767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8048__B _3059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6347__I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_61 io_oeb[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__7774__A2 _2903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8971__A1 _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6577__A3 _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_as2650_72 io_oeb[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_3398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_83 io_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5785__A1 _4228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_94 io_oeb[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_109_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9246__CLK clknet_leaf_62_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8487__B1 _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4760__A2 _4225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7641__I _2520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7462__A1 _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7830_ as2650.pc\[10\] _1586_ _2959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_58_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7761_ _2788_ _2891_ _2843_ _2892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4973_ _4154_ _4552_ _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6712_ as2650.stack\[0\]\[11\] _1927_ _1930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7692_ _2573_ _2824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_75_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7517__A2 _2532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8714__A1 _3763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6643_ _1838_ _1849_ _1872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5528__A1 _4375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7816__I net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8190__A2 _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9362_ _0255_ clknet_leaf_69_wb_clk_i as2650.r123\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6574_ _4519_ _1783_ _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8313_ _2437_ _3415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5525_ _0829_ _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_9293_ _0186_ clknet_leaf_20_wb_clk_i net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8244_ _3089_ _2438_ _3344_ _3346_ _3347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_69_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5456_ _0760_ _0761_ _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8175_ _2336_ _0885_ _1462_ _3279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5700__A1 as2650.stack\[6\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7551__I _1513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5387_ _0505_ _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7126_ _2215_ _2175_ _2291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7453__A1 _2584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6256__A2 _1513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7057_ as2650.r123_2\[3\]\[6\] _2241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9119__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6008_ _4214_ _4250_ _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7205__A1 _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6008__A2 _4250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7756__A2 _2886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8953__A1 _3995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5767__A1 _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7959_ _2149_ _3081_ _3083_ _3084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5020__B _4454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5519__A1 _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4990__A2 _4385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8181__A2 _3163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7461__I _2564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6247__A2 _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7995__A2 _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8795__I1 _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6955__B1 _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6026__B _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4981__A2 _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8172__A2 _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9056__C _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7380__B1 _2516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5310_ _4426_ _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6290_ _1546_ _1547_ _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5369__S0 _4196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9072__B _4105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5241_ as2650.holding_reg\[4\] _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5172_ _0480_ _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6238__A2 _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput2 io_in[11] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8931_ _3981_ _3982_ _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8416__B _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8862_ _2285_ _3931_ _3932_ as2650.stack\[7\]\[1\] _3933_ _3934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_37_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8935__A1 _4272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7813_ _1565_ _2943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5749__A1 _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8793_ _2635_ _1537_ _1450_ _3876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7744_ _1616_ _0829_ _2875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4956_ _4397_ _4535_ _4536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7675_ _0683_ _0697_ _2808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4972__A2 _4242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4887_ _4467_ _4458_ _4468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_138_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8163__A2 _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6450__I _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6626_ _1838_ _1849_ _1855_ _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_14_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6174__A1 _4303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7910__A2 _2504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9345_ _0238_ clknet_leaf_52_wb_clk_i as2650.stack\[6\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6557_ _1756_ _1766_ _1788_ _1789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_14_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5921__A1 _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5066__I _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5508_ as2650.holding_reg\[7\] _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9276_ _0169_ clknet_3_2_0_wb_clk_i as2650.addr_buff\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6488_ _4405_ _1723_ _1724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_134_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7674__A1 _2800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8227_ _3287_ _3331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5439_ _0599_ _0744_ _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8158_ net4 _3263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_126_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6229__A2 _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7109_ as2650.r123\[3\]\[7\] _2276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8089_ _3193_ _3197_ _3198_ _3200_ _2624_ _3201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_101_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7977__A2 _3087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5988__A1 _4215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4660__A1 _4237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8926__A1 _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6165__A1 as2650.stack\[4\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4715__A2 _4198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9103__A1 as2650.psu\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7665__A1 _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7124__C _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8090__A1 _3178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5979__A1 _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8393__A2 _3457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4810_ _4390_ _4391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7794__C _2923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5790_ _1070_ _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_56_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4741_ _4321_ _4311_ _4322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7366__I _2504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7460_ _2560_ _2596_ _2597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4672_ _4251_ as2650.cycle\[2\] _4252_ _4253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_135_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6411_ _1659_ _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7391_ _1260_ _0872_ _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9130_ _0023_ clknet_leaf_58_wb_clk_i as2650.stack\[5\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6342_ _0835_ _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_116_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7656__A1 _2785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9061_ _1575_ _4010_ _4096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7315__B _2453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6273_ _1530_ _1273_ _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8012_ _3131_ _0192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5224_ _0526_ _0530_ _0531_ _0532_ _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_29_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7408__A1 _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5155_ _0463_ _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_99_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7959__A2 _3081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8081__A1 _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8081__B2 _3154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5086_ _0395_ _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6631__A2 _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8914_ _3968_ _3970_ _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8908__A1 _4414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8845_ _2265_ _3904_ _3906_ as2650.stack\[6\]\[6\] _3910_ _3920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_38_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8384__A2 _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_77_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6395__A1 _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8776_ _2399_ _0639_ _2514_ _3860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5988_ _4215_ _4223_ _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7727_ _2854_ _2856_ _2857_ _2858_ _2859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_40_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4939_ as2650.r0\[2\] _4519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7276__I _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6147__A1 _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7658_ _2778_ _2542_ _2499_ _2791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7895__A1 _2998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6609_ _4382_ _1811_ _1839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7589_ _2191_ _2684_ _2723_ _2681_ _2724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_105_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_opt_1_0_wb_clk_i clknet_3_6_0_wb_clk_i clknet_opt_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_9328_ _0221_ clknet_3_7_0_wb_clk_i as2650.pc\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_21_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5370__A2 _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7647__A1 _2778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9259_ _0152_ clknet_leaf_55_wb_clk_i as2650.stack\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4881__A1 as2650.stack\[2\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8056__B _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6355__I _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6622__A2 _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8375__A2 _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9318__D _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8127__A2 _3236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8011__S _3130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8835__B1 _3909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5113__A2 _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6310__A1 _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8063__A1 _2618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6265__I _4428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6613__A2 _4284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6960_ _2139_ _1657_ _2166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_81_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5911_ _0668_ _1060_ _1187_ _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6891_ _1794_ _2100_ _2101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8366__A2 _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8630_ _3329_ _3706_ _3721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5842_ _1093_ _1055_ _1122_ _0031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8561_ _2527_ _3652_ _3654_ _2160_ _3655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_37_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5773_ _1054_ _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5609__I _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7512_ _2384_ _2648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4724_ _4283_ _4305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8492_ _3317_ _3563_ _3580_ _3582_ _3588_ _2391_ _3589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
X_7443_ _2517_ _2580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4655_ _4173_ as2650.cycle\[0\] _4236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7374_ _2492_ _2513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5352__A2 _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4586_ _4163_ _4166_ _4167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_11_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7629__A1 _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9113_ _0006_ clknet_leaf_67_wb_clk_i as2650.r123\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6325_ _1581_ _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_66_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5344__I _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9044_ _0299_ _0319_ _4343_ _4080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6256_ _0814_ _1513_ _1266_ _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_107_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5207_ _4220_ _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6187_ _0408_ _0445_ _0543_ _0641_ _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_69_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4863__A1 _4443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8054__A1 _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5138_ _0393_ _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7801__A1 _2926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6604__A2 _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5069_ _4399_ _0378_ _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6368__A1 _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8828_ _3903_ _3908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8759_ _1235_ _3844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8109__A2 _3212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5591__A2 _4208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6540__B2 _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5254__I _4338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8832__A3 _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8596__A2 _3687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4606__A1 as2650.ins_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4909__A2 _4489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7859__A1 _2369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7644__I _2776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8520__A2 _3596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7323__A3 _2461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5164__I _4279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6110_ _0337_ _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7090_ _2265_ _2247_ _2250_ as2650.stack\[1\]\[6\] _2254_ _2266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_112_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6041_ _4235_ _4241_ _1313_ _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4845__A1 _4420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_47_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_47_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_67_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7992_ _1550_ _1442_ _3114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6598__A1 _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9152__CLK clknet_leaf_16_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6943_ _0873_ _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8339__A2 _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6874_ _1970_ _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8613_ _1002_ _0995_ _3663_ _3704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7011__A2 _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5825_ _0301_ _4534_ _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5022__A1 as2650.stack\[0\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8544_ _3638_ _3639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5756_ _4189_ _1037_ _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4707_ _4285_ _4140_ _4286_ _4287_ _4288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_136_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8475_ _2925_ _3163_ _3156_ _3572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7554__I net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5275__S _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5687_ _0971_ _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8511__A2 _4370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7426_ _1341_ _2564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6522__A1 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5325__A2 _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4638_ _4215_ _4218_ _4219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_89_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7357_ _2492_ _2495_ _2496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5074__I _4503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4569_ _4149_ _4150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_144_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8275__A1 _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6308_ _1565_ _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_81_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7288_ _1471_ _1501_ _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5089__A1 as2650.holding_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8814__A3 _3895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9027_ _1475_ _2447_ _4060_ _4063_ _4064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_134_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6239_ _4255_ _1497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8578__A2 _3665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7250__A2 _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5261__A1 _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7305__A3 _2443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6513__A1 _4284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9331__D _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4827__A1 _4154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9175__CLK clknet_leaf_60_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8228__C _3331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8569__A2 _3621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5252__A1 _4488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9059__C _3742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5004__A1 _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5610_ _0902_ _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6590_ _1801_ _1804_ _1820_ _1821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__5555__A2 _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5541_ _0296_ _0821_ _0845_ _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7374__I _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8260_ as2650.stack\[2\]\[1\] _1637_ _3363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5307__A2 _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6504__A1 as2650.r123_2\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5472_ as2650.stack\[0\]\[14\] _4465_ _4469_ as2650.stack\[1\]\[14\] _0778_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_144_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6504__B2 _1738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7211_ _2334_ _2358_ _2360_ _0162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8191_ _1544_ _2487_ _3294_ _3295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7142_ _2302_ _2281_ _2283_ as2650.stack\[3\]\[5\] _2278_ _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_113_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7073_ _2243_ _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6024_ as2650.psu\[5\] _1292_ _1295_ _1297_ _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7480__A2 _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7042__C _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7232__A2 _2363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7975_ _3088_ _3098_ _3099_ _2923_ _3100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_82_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7549__I _2517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5243__A1 _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8980__A2 _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6926_ _0791_ _2109_ _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6991__A1 _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6857_ _2037_ _2040_ _2067_ _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xfanout46 net48 net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__8732__A2 _3766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5808_ _1089_ _0969_ _4492_ _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6788_ _4366_ _1763_ _2001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6743__A1 _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8527_ _0964_ _3594_ _3622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5739_ _0985_ _1022_ _1026_ _0024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8496__A1 _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8458_ _4477_ _3553_ _3554_ _3555_ _3556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_136_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7409_ _2530_ _1619_ _2499_ _2546_ _2547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_8389_ _3481_ _3488_ _3489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9198__CLK clknet_leaf_46_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8248__A1 _3048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8248__B2 _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8799__A2 _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5532__I _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8420__A1 as2650.stack\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8064__B _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_62 io_oeb[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_3399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8971__A2 _2509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_73 io_oeb[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_84 io_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5785__A2 _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6982__A1 _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_as2650_95 io_oeb[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6734__A1 _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5707__I _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4611__I _4183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8487__B2 as2650.stack\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7922__I _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8239__A1 _2777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8753__I _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8411__A1 _2736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7369__I _2507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7760_ _2783_ _2842_ _2891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4972_ _4551_ _4242_ _4246_ _4552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_63_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6711_ _1666_ _1924_ _1929_ _0093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7691_ _2774_ _2822_ _2823_ _0179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8714__A2 _3788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6642_ _1838_ _1849_ _1871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_123_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9361_ _0254_ clknet_leaf_74_wb_clk_i as2650.r123\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6573_ _1782_ _1802_ _1803_ _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5617__I as2650.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8312_ _3070_ _3407_ _3413_ _3414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8478__A1 _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5524_ _4375_ _0487_ _0822_ _0571_ _0825_ _4358_ _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
X_9292_ _0185_ clknet_leaf_31_wb_clk_i net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9340__CLK clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8243_ _4531_ _3345_ _3346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5455_ _4218_ _0638_ _0664_ _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_105_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_62_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_62_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_8174_ _2631_ _3274_ _3275_ _3277_ _3278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__5700__A2 _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5386_ _4515_ _0681_ _0692_ _4538_ _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__8149__B _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7125_ _1382_ _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7056_ _2240_ _0127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6256__A3 _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5464__A1 _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6007_ _4430_ _1280_ _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5464__B2 _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8402__A1 _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7205__A2 _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7279__I _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8953__A2 _2076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7958_ _1482_ _1293_ _2160_ _3082_ _3083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6964__A1 _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6909_ as2650.r123_2\[2\]\[5\] _2019_ _2117_ _1980_ _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7889_ _2974_ _3014_ _3015_ _2961_ _3016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_23_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8181__A3 _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5262__I _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6247__A3 _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5455__A1 _4218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9213__CLK clknet_leaf_56_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6955__A1 _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5758__A2 _4198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6955__B2 _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_46_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9363__CLK clknet_leaf_69_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8172__A3 _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7380__A1 _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5369__S1 _4148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5240_ _0414_ _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6268__I _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5171_ _4518_ _4523_ _0365_ _0368_ _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_68_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8632__A1 _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8930_ _0775_ _3958_ _3982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput3 io_in[12] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5900__I as2650.r123_2\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7199__A1 _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8861_ _3923_ _3933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8935__A2 _1612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7812_ _2465_ _2942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8792_ _3804_ _0749_ _3874_ _3875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6946__A1 _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7743_ _2870_ _2873_ _2874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4955_ _4387_ _4534_ _4535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_33_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8699__A1 _3143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7674_ _2800_ _0697_ _2807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_127_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4886_ as2650.psu\[0\] _4467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5057__S0 _4139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4972__A3 _4246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6625_ _1850_ _1852_ _1854_ _1855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_53_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7371__A1 _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6174__A2 _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7990__C _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6556_ _0492_ _1722_ _1750_ _1788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_20_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9344_ _0237_ clknet_leaf_37_wb_clk_i as2650.stack\[6\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5382__B1 _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5507_ _0313_ _0811_ _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9275_ _0168_ clknet_leaf_11_wb_clk_i as2650.addr_buff\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6487_ _1722_ _1723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8226_ _3316_ _3328_ _3329_ _3330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7674__A2 _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5438_ _0502_ _0588_ _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8157_ as2650.psu\[7\] _3262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_82_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5369_ as2650.r123\[1\]\[6\] as2650.r123\[0\]\[6\] as2650.r123_2\[1\]\[6\] as2650.r123_2\[0\]\[6\]
+ _4196_ _4148_ _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_59_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7108_ _2275_ _0144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6229__A3 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8088_ _2383_ _3192_ _3169_ _3199_ _3200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_43_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7511__B _2646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7039_ _2193_ _2211_ _2231_ _0119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_142_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5988__A2 _4223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4660__A2 _4240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8926__A2 _3969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9386__CLK clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_output15_I net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8342__B _3442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7362__A1 _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6165__A2 _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5257__I _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7665__A2 _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8862__A1 _2285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5676__A1 _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5428__A1 _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7421__B _2554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8090__A2 _3192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_2_wb_clk_i_I clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5876__B _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4740_ _4320_ as2650.carry _4321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9067__C _4097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8145__A3 as2650.cycle\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4671_ as2650.cycle\[1\] as2650.cycle\[0\] _4252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6410_ _1658_ _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9109__CLK clknet_leaf_68_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7390_ _2525_ _2527_ _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6341_ as2650.psl\[1\] _1104_ _1588_ _1525_ _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__9083__B _3619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7382__I _2464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9060_ _3106_ _1046_ _1244_ _2631_ _4095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__7656__A2 _2788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6272_ _0751_ _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_66_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8011_ _3129_ _0413_ _3130_ _3131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__9259__CLK clknet_leaf_55_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5223_ as2650.stack\[7\]\[11\] _4478_ _0527_ as2650.stack\[6\]\[11\] _0329_ _0532_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_102_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7408__A2 _2545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8605__A1 _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5154_ _0462_ _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4890__A2 _4466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8081__A2 _3192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5085_ _0393_ _0394_ _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_96_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6092__A1 _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8913_ _0323_ _3969_ _3970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8908__A2 _3959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9030__A1 _3827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8844_ _0938_ _3902_ _3919_ _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_53_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7592__A1 _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8775_ _3804_ _0668_ _3858_ _3859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5987_ _4369_ _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6395__A2 _1643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7726_ net54 _2505_ _2688_ _2542_ _2858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4938_ _4297_ _4517_ _4518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7657_ _2784_ _2789_ _2790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7344__A1 _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4869_ _4449_ _4450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6608_ _4294_ _1812_ _1808_ _1838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_7588_ _2685_ _2702_ _2722_ _2723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7895__A2 _2871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9327_ _0220_ clknet_3_7_0_wb_clk_i as2650.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6539_ _1771_ _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__9097__A1 _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8844__A1 _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9258_ _0151_ clknet_leaf_56_wb_clk_i as2650.stack\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5658__A1 _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8209_ _3293_ _3308_ _3312_ _3313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_133_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9189_ _0082_ clknet_leaf_65_wb_clk_i as2650.r123_2\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4881__A2 _4461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8056__C _2482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5830__A1 _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8851__I _3923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9021__A1 _4491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6371__I _1480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9088__A1 _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9334__D _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8835__A1 _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5651__S _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8063__A2 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6074__A1 _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4624__A2 _4204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5910_ _1136_ _1185_ _1186_ _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__9012__A1 _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6890_ _2097_ _2099_ _2100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_62_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5841_ _1056_ _1116_ _1121_ _1054_ _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_62_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7574__A1 _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8560_ _2365_ _2776_ _3653_ _3654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5772_ _1053_ _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7511_ _2643_ _2644_ _2646_ _2647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4723_ _4283_ _4289_ _4304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
X_8491_ _3583_ _3584_ _3587_ _3588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8710__B _3797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7442_ _2520_ _2579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4654_ _4234_ _4235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5888__A1 _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7373_ _2498_ _2500_ _2502_ _2511_ _2512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_128_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9079__A1 _4365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4585_ _4165_ _4166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6324_ _1580_ _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_9112_ _0005_ clknet_leaf_68_wb_clk_i as2650.r123\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7629__A2 _2762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8826__A1 _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9043_ _0299_ _0320_ _4079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6255_ _1471_ _1513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_118_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5206_ _4389_ _0505_ _0514_ _4221_ _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_48_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6186_ _4258_ _1440_ _1441_ _1443_ _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_57_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4863__A2 _4426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5137_ _0395_ _0445_ _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8054__A2 _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6065__A1 _4238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7996__B _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7801__A2 _2928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5068_ _4525_ _0377_ _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_44_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9003__A1 _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8827_ _0848_ _3902_ _3907_ _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_77_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7565__A1 _2687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6368__A2 _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4704__I _4284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8758_ _0619_ _3488_ _3843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_139_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5040__A2 _4509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7709_ _2720_ _2840_ _2818_ _2841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7317__A1 _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8689_ _3768_ _3776_ _3777_ _3778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6540__A2 _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8817__A1 _3837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6366__I _4219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5270__I _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5803__A1 _4472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7556__A1 _2687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7308__A1 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6969__C _2173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5319__B1 _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4790__A1 _4369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5873__C _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5445__I _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5185__I3 as2650.r123_2\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8808__A1 _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7660__I _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6040_ _1308_ _1312_ _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input6_I io_in[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4845__A2 _4422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7991_ _4406_ _1524_ _3113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6942_ _0957_ _2148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_16_wb_clk_i clknet_3_3_0_wb_clk_i clknet_leaf_16_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_35_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7547__A1 _2643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6873_ _0586_ _2005_ _2083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8612_ _2415_ _3703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5824_ _1072_ _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5022__A2 _4465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8543_ _3257_ _3624_ _3630_ _2549_ _2928_ _3638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_33_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5755_ _4143_ _1036_ _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4706_ as2650.r123\[1\]\[0\] as2650.r123\[0\]\[0\] as2650.r123_2\[1\]\[0\] as2650.r123_2\[0\]\[0\]
+ as2650.ins_reg\[0\] _4146_ _4287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_8474_ _2203_ _3570_ _3571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5686_ _4415_ _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7425_ _2473_ _2562_ _2563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4637_ _4217_ _4218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5355__I _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7356_ _2494_ _2495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4568_ _4148_ _4149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6307_ _4203_ _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8275__A2 _3377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7287_ _2422_ _2425_ _2426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5089__A2 _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6238_ _1316_ _1275_ _1357_ _1496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_9026_ _1463_ _4061_ _4062_ _4063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_57_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6169_ _4344_ _0321_ _0422_ _0476_ _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_58_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7786__A1 _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7250__A3 _1702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8334__C _3434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5261__A2 _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7538__A1 _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6210__A1 _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7710__A1 as2650.pc\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6029__A1 _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6029__C _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7777__A1 _2889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5252__A2 _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6201__A1 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5555__A3 _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5540_ _0700_ _0828_ _0831_ _0844_ _0295_ _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_34_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5471_ as2650.stack\[4\]\[14\] _4481_ _0430_ as2650.stack\[5\]\[14\] _0329_ _0777_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_69_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6504__A2 _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7701__A1 _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7210_ _1691_ _2359_ _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8190_ _2144_ _1605_ _3294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7604__B _2737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7141_ _2196_ _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8257__A2 _4474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5903__I _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7072_ _2249_ _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6023_ _1291_ _1296_ _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7974_ net51 _3090_ _2155_ _3099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5243__A2 _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6440__A1 _4223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6925_ _2122_ _2128_ _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_74_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8980__A3 _4016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6856_ _4367_ _1764_ _2041_ _2067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xfanout47 net48 net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_126_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5807_ _0294_ _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7940__A1 _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6787_ _4366_ _1749_ _1764_ _0672_ _2000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6743__A2 _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8526_ _3288_ _3621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4754__A1 _4332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5738_ as2650.stack\[5\]\[9\] _1025_ _1026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8496__A2 _3289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8457_ as2650.stack\[4\]\[6\] _1904_ _1656_ as2650.stack\[5\]\[6\] _4476_ _3555_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5669_ _0964_ _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7408_ _2542_ _2545_ _2546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8388_ _3482_ _3483_ _3484_ _3487_ _3488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_137_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7339_ _2467_ _2471_ _2475_ _2477_ _2478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_116_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9009_ _4039_ _4046_ _4047_ _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_3301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7759__A1 as2650.pc\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8420__A2 _2215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_63 io_oeb[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_3389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8971__A3 _3048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_36_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_as2650_74 io_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8708__B1 _4435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xwrapped_as2650_85 io_oeb[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_2677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6982__A2 _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4993__A1 as2650.holding_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7475__I _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6734__A2 _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4745__A1 _4303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5209__B _4545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8487__A2 _1905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9142__CLK clknet_leaf_67_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5170__A1 _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8239__C _3089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9292__CLK clknet_leaf_31_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_75_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6670__A1 _1795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8411__A2 _2756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5225__A2 _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4971_ _4550_ _4551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_92_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6710_ as2650.stack\[0\]\[10\] _1927_ _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4984__A1 _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7690_ _2778_ _2771_ _2772_ _2823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8175__A1 _2336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9086__B as2650.psl\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6641_ _1850_ _1868_ _1869_ _1870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4802__I _4382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4736__A1 as2650.psl\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9360_ _0253_ clknet_leaf_59_wb_clk_i as2650.stack\[7\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6572_ _1785_ _1786_ _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_125_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8311_ _3093_ _3412_ _3413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5523_ _0827_ _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_9291_ _0184_ clknet_leaf_31_wb_clk_i net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8478__A2 _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6489__A1 _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8242_ _2533_ _3345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5454_ _4533_ _0589_ _0574_ _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_117_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5161__A1 _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5385_ _0685_ _4532_ _0691_ _4378_ _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_8173_ _2428_ _3276_ _3277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7124_ _2285_ _2286_ _2287_ as2650.stack\[3\]\[1\] _2288_ _2289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_141_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7055_ as2650.r123_2\[3\]\[5\] _2240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6661__A1 _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6006_ _1278_ _0418_ _1279_ _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__5464__A2 _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_31_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_31_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_74_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8402__A2 _2539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6413__A1 as2650.stack\[2\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5301__C _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7957_ _2493_ _3082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6908_ _2103_ _2105_ _2116_ _2117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_7888_ as2650.pc\[11\] _0988_ _2825_ _3015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6839_ _2023_ _2046_ _2050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7913__A1 _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6716__A2 _1923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8181__A4 _3065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4727__A1 _4305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9165__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8509_ _2996_ _3595_ _3605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_87_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5527__I0 _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9162__D _0055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8854__I _3926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6247__A4 _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6652__A1 as2650.r0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5455__A2 _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6955__A2 _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5758__A3 _4151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8522__C _3420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7904__A1 _2963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9337__D _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5718__I _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4622__I _4202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7380__A2 _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7933__I _3058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5143__A1 _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5453__I _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6340__B1 _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6891__A1 _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5170_ _0477_ _0478_ _0352_ _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_96_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8632__A2 _3377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput4 io_in[13] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_42_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8860_ _3928_ _3932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7199__A2 _2348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7811_ _0979_ _2684_ _2939_ _2940_ _2941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8791_ _2565_ _0771_ _3874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7742_ _2334_ _2872_ _2873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4957__A1 _4531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8148__A1 _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9188__CLK clknet_leaf_69_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4954_ _4217_ _4533_ _4333_ _4534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_51_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7673_ _1587_ _0770_ _2806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_33_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8699__A2 _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4885_ _4465_ _4466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5057__S1 _4516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4709__A1 _4190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6624_ _1853_ _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7371__A2 _2509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9343_ _0236_ clknet_leaf_38_wb_clk_i as2650.stack\[6\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5382__A1 _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6555_ _1782_ _1785_ _1786_ _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_119_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5382__B2 _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5506_ _4336_ _0810_ _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9274_ _0167_ clknet_leaf_11_wb_clk_i as2650.addr_buff\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8320__A1 _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6486_ _1721_ _1722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8225_ _3290_ _3329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6459__I _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5134__A1 as2650.holding_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5437_ _0741_ _0742_ _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5363__I _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8156_ _3208_ _1329_ _3229_ _3261_ _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5368_ _4369_ _0674_ _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7107_ as2650.r123\[3\]\[6\] _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8674__I _3757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5299_ _4364_ _0372_ _0606_ _4362_ _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_8087_ _3170_ _3199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6229__A4 _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7038_ _2197_ _2214_ _2217_ as2650.stack\[4\]\[5\] _2210_ _2231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_28_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8387__A1 as2650.stack\[7\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6127__C _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_28_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8989_ _0849_ _0426_ _4029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8342__C _3058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7362__A2 _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7753__I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8311__A1 _3093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7114__A2 _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5125__A1 _4477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8862__A2 _3931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6873__A1 _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5206__C _4221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8075__B1 _3185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5428__A2 _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8378__A1 _3472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9330__CLK clknet_leaf_80_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8025__S _3130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5448__I _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4670_ as2650.cycle\[3\] _4251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8759__I _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6561__B1 _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6340_ as2650.overflow _0375_ _1594_ _4320_ _1596_ _1597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_115_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6271_ _1525_ _1526_ _1527_ _1528_ _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6279__I _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5183__I _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5222_ as2650.stack\[4\]\[11\] _0429_ _0430_ as2650.stack\[5\]\[11\] _0531_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8010_ _3119_ _3130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_130_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5153_ _0365_ _0368_ _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_96_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6616__A1 as2650.r0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5419__A2 _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5084_ _4278_ _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6092__A2 _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8912_ _3958_ _3969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8369__A1 _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8843_ _2302_ _3904_ _3906_ as2650.stack\[6\]\[5\] _3901_ _3919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_20_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9030__A2 _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7041__A1 _2200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8774_ _2598_ _0698_ _3858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5986_ _4393_ _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7592__A2 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7725_ _2648_ _2840_ _2857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4937_ as2650.r123\[2\]\[2\] as2650.r123_2\[2\]\[2\] _4516_ _4517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_123_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7656_ _2785_ _2788_ _2789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4868_ as2650.psu\[0\] as2650.psu\[1\] _4449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8541__A1 _3572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7344__A2 _2482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8541__B2 _3395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6607_ _1814_ _1819_ _1837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8669__I _3757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7587_ _1337_ _2715_ _2718_ _2719_ _2721_ _2722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__7895__A3 _2868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4799_ as2650.r123\[2\]\[1\] as2650.r123_2\[2\]\[1\] _4379_ _4380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_107_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9326_ _0219_ clknet_3_6_0_wb_clk_i as2650.pc\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6538_ _1767_ _1770_ _1771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_14_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__9097__A2 _3144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5107__A1 _4315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9203__CLK clknet_leaf_47_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9257_ _0150_ clknet_leaf_55_wb_clk_i as2650.stack\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6469_ _4160_ _1688_ _1698_ _1706_ _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_121_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8208_ _0864_ _2854_ _3058_ _3311_ _3312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5658__A2 _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9188_ _0081_ clknet_leaf_69_wb_clk_i as2650.r123_2\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8139_ _3243_ _3244_ _3247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5821__I _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9353__CLK clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8072__A3 _3184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7280__A1 _4199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9021__A2 _3268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8780__A1 _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8532__A1 _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7335__A2 _4361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8800__C _2630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5897__A2 _1174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9088__A2 _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8835__A2 _3908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6074__A2 _4237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7271__A1 _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5840_ _0344_ _1117_ _1120_ _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_61_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7574__A2 _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5585__A1 _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5771_ _4437_ _1035_ _1052_ _4438_ _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__5178__I _4359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7510_ _1684_ _2645_ _2646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4722_ _4290_ _4293_ _4302_ _4303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_37_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8490_ as2650.stack\[6\]\[7\] _1639_ _4476_ _3586_ _3587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_30_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7441_ _2521_ _2575_ _2576_ _2578_ _0174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_30_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5337__A1 _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4653_ as2650.cycle\[7\] _4234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__9226__CLK clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4810__I _4390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7372_ _2418_ _2505_ _2508_ _1551_ _2510_ _2511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4584_ as2650.cycle\[3\] _4164_ _4165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_9111_ _0004_ clknet_leaf_68_wb_clk_i as2650.r123\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6323_ _0595_ _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_89_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9376__CLK clknet_leaf_74_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6837__B2 _1980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9042_ _1691_ _4056_ _4070_ _4078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6254_ _1488_ _1491_ _1506_ _1511_ _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_131_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5205_ _0508_ _4399_ _0513_ _4230_ _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5641__I _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6185_ _1442_ _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5136_ _0444_ _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8054__A3 _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7262__A1 _4323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6065__A2 _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5067_ _4218_ _4507_ _4510_ _4533_ _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7996__C _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9003__A2 _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6472__I _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8826_ _2146_ _3904_ _3906_ as2650.stack\[6\]\[0\] _3901_ _3907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_77_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7565__A2 _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5576__A1 _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8757_ _3838_ _0570_ _3184_ _3840_ _3841_ _3842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5969_ _4137_ _1242_ _4425_ _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7708_ _2838_ _2839_ _2840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_138_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8688_ _4219_ _3777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8514__A1 _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7317__A2 _2430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7517__B _2652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7639_ _2757_ _2771_ _2772_ _2773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5816__I _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9309_ _0202_ clknet_leaf_16_wb_clk_i as2650.cycle\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_107_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8817__A2 _3897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5803__A2 _4484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6382__I _1637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7556__A2 _2690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9249__CLK clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7308__A2 _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5319__A1 as2650.stack\[0\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4790__A2 _4370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5319__B2 as2650.stack\[1\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4630__I _4210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8808__A2 _3588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7492__A1 _2579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4845__A3 _4425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7990_ _3107_ _3110_ _3111_ _3112_ _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_93_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5255__B1 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8992__A1 _2794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6941_ _2146_ _2147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_35_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6292__I _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6872_ _2060_ _2080_ _2081_ _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_39_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7547__A2 _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8744__A1 _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8611_ _3035_ _3374_ _3701_ _3702_ _2415_ _0220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__8744__B2 _4434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5823_ _4529_ _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_8542_ _3625_ _3627_ _3636_ _3637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5754_ _4248_ _4151_ _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_56_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_56_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_31_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4705_ _4138_ _4135_ _4286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8473_ _0945_ _2195_ _2187_ _3427_ _3570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_72_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5685_ _0967_ _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7424_ _4529_ _4513_ _2561_ _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_120_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4636_ _4182_ _4216_ _4217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7355_ _2493_ _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4567_ _4147_ _4148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6306_ _1449_ _1461_ _1563_ _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_85_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7286_ _2419_ _2424_ _4418_ _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8168__B _3229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9025_ _2395_ _1264_ _4062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6237_ _1323_ _1493_ _1494_ _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_83_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6168_ _1016_ _1418_ _1426_ _0053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_58_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7235__A1 _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5119_ _4465_ _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_79_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6099_ _1334_ _1353_ _1366_ _1371_ _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_100_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_17_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8983__A1 _3844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5797__A1 _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_26_wb_clk_i_I clknet_opt_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8035__I0 _3149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_3_3_0_wb_clk_i clknet_0_wb_clk_i clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_41_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6135__C _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7538__A2 _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8735__A1 _3703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8809_ _1611_ _3793_ _3891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6210__A2 _4431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5546__I _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7710__A2 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6578__S _4144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7474__A1 _2609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6377__I _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5281__I _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_65_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8806__B _3887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6029__A2 _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8423__B1 _3386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8974__A1 _3045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5788__A1 _4395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5230__B _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7001__I _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8726__A1 _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5470_ as2650.stack\[7\]\[14\] _0326_ _0527_ as2650.stack\[6\]\[14\] _0776_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_129_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7701__A2 _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5712__A1 _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7140_ _2186_ _2279_ _2301_ _0150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7604__C _2662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6287__I _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5191__I _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7071_ _2246_ _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6022_ _4199_ _1264_ _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_140_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8965__A1 _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7973_ _3092_ _3097_ _3098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6924_ _2107_ _2114_ _2127_ _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_70_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6440__A2 _1681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8980__A4 _4019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6855_ _2062_ _2065_ _2066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_23_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout48 net49 net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_11_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5806_ _1087_ _1036_ _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6786_ _1964_ _1997_ _1998_ _1999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7940__A2 _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8525_ _2911_ _3620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5737_ _1020_ _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4754__A2 _4334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8456_ as2650.stack\[7\]\[6\] _3366_ _3386_ as2650.stack\[6\]\[6\] _3554_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_5668_ as2650.pc\[8\] _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_11_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7407_ _2543_ _2544_ _2545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4619_ as2650.halted _4200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8677__I _3765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8387_ as2650.stack\[7\]\[4\] _1920_ _3486_ _3487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5599_ _0902_ _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7338_ _2476_ _2477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7456__A1 _4511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5315__B _4454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7269_ _1260_ _1248_ _2409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_133_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9008_ _4463_ _4039_ _1634_ _4047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_77_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5219__B1 _4469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8956__A1 _3976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4690__A1 _4213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output38_I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_64 io_oeb[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__8971__A4 _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_75 io_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8708__A1 _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_86 io_oeb[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_109_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4993__A2 _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6195__A1 _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5942__A1 _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4745__A2 _4310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7705__B _2836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_1_wb_clk_i clknet_3_0_0_wb_clk_i clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_126_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5170__A2 _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8644__B1 _3733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6670__A2 _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4681__A1 _4248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8255__C _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8947__A1 _3995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4970_ _4232_ _4550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_36_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4984__A2 _4261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8175__A2 _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6640_ _1852_ _1854_ _1869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6186__A1 _4258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6571_ _1785_ _1786_ _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4736__A2 _4316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8310_ _3082_ _3381_ _3409_ _2645_ _3411_ _3412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_118_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5522_ _0823_ _0826_ _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9290_ _0183_ clknet_leaf_28_wb_clk_i net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7686__A1 _2613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8241_ _2362_ _3181_ _3344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6489__A2 _4152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7686__B2 _2818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5453_ _0758_ _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8172_ _0853_ _1248_ _2427_ _3276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_114_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5161__A2 _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5384_ _0598_ _0690_ _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7438__A1 _2530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7123_ _2277_ _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7054_ _2239_ _0126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8446__B _3543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7350__B _2483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6005_ _1262_ _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8938__A1 _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6413__A2 _1661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7956_ _1617_ _2352_ _3081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_71_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_71_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_42_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6907_ _2115_ _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_42_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7887_ _3013_ _3014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_126_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4975__A2 _4513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6838_ _1139_ _1938_ _2049_ _0100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5924__A1 _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4727__A2 _4306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6769_ _1116_ _1940_ _1942_ as2650.r123_2\[2\]\[1\] _1982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_137_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8508_ _2334_ _2755_ _1509_ _3603_ _3604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_104_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8439_ _0758_ _0674_ _3537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_137_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6652__A2 _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5455__A3 _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8075__C _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9051__B1 _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7601__A1 _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6955__A3 _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6168__A1 _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4718__A2 _4281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7668__A1 _2800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5734__I _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5143__A2 _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6340__B2 _4320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6891__A2 _2100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8093__A1 _3186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6643__A2 _1849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput5 io_in[33] net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7810_ _1327_ _2940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8790_ _3837_ _3872_ _3873_ _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_91_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7741_ _2871_ _2869_ _2872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9097__B _4121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4953_ _4249_ _4258_ _4533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__8148__A2 _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7672_ _1559_ _2553_ _2467_ _2804_ _2805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_36_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4884_ _4464_ _4465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6623_ _0671_ _1721_ _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5906__A1 _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9342_ _0235_ clknet_leaf_38_wb_clk_i as2650.stack\[6\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6554_ _0499_ _1721_ _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5382__A2 _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7659__A1 _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5505_ _0550_ _4376_ _0809_ _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_9273_ _0166_ clknet_leaf_12_wb_clk_i as2650.addr_buff\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6485_ _1720_ _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8320__A2 _3377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8224_ _0864_ _3317_ _3326_ _3327_ _3328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_133_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5436_ _0590_ _0686_ _0678_ _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5134__A2 _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8155_ _1570_ _3257_ _3258_ _3260_ _3207_ _3261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA_clkbuf_3_1_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5367_ as2650.r123\[2\]\[6\] as2650.r123_2\[2\]\[6\] _0493_ _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_47_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8084__A1 _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7106_ _2274_ _0143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8086_ _2399_ _3167_ _3198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8623__A3 _3713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8176__B _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5298_ _4378_ _0593_ _0605_ _4222_ _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_87_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6634__A2 _1858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7037_ _2186_ _2211_ _2230_ _0118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4645__A1 _4192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8387__A2 _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9132__CLK clknet_leaf_56_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8988_ _2634_ _3266_ _4028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7939_ net49 _3056_ _3064_ _2578_ _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5070__A1 _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5819__I _4334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7898__A1 _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9282__CLK clknet_leaf_26_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6570__A1 _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7255__B _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8698__I0 _4513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8847__B1 _3909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5676__A3 _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8075__A1 _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8075__B2 _3187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8105__I _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7889__A1 _2974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8550__A2 as2650.pc\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8838__B1 _3909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6270_ _1239_ _0759_ _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5221_ as2650.stack\[0\]\[11\] _0429_ _0527_ as2650.stack\[2\]\[11\] _0529_ _0530_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_69_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8066__A1 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8708__C _3777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5152_ as2650.holding_reg\[3\] _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6295__I _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6616__A2 _1730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4808__I _4229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5083_ _4312_ _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8911_ _3966_ _1738_ _3967_ as2650.r123\[1\]\[1\] _3968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_49_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8369__A2 _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8842_ _0932_ _3902_ _3918_ _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_64_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8773_ _3837_ _3855_ _3857_ _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5985_ _1249_ _1258_ _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7724_ _2855_ _2856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4936_ _4147_ _4516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_36_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7655_ _2786_ _2787_ _2788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_21_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4867_ as2650.psu\[2\] _4448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7854__I net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8541__A2 _3624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6606_ _1815_ _1834_ _1835_ _1836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7586_ _2720_ _2691_ _2570_ _2721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6552__A1 _4382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6552__B2 _4284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4798_ _4145_ _4379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7895__A4 _3021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9325_ _0218_ clknet_leaf_30_wb_clk_i as2650.pc\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6537_ _1768_ _1769_ _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5374__I _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9256_ _0149_ clknet_leaf_44_wb_clk_i as2650.stack\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6304__A1 _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6468_ _1559_ _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8207_ _2382_ _3310_ _3311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5419_ _0649_ _0720_ _0722_ _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_9187_ _0080_ clknet_leaf_65_wb_clk_i as2650.r123_2\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6399_ _1006_ _1644_ _1650_ _0060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_121_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4866__A1 _4441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8138_ _3243_ _3244_ _3246_ _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_47_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8069_ _1272_ _3181_ _3182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9006__B1 _4044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7280__A2 _4544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5291__A1 _4508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6933__I _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5043__A1 _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8780__A2 _3793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8517__C1 _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6791__A1 _4519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5346__A2 _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5284__I _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9088__A3 _4062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8296__A1 _3382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9178__CLK clknet_leaf_73_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8048__A1 _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7004__I as2650.pc\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7271__A2 _1513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_opt_1_0_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5034__A1 _4494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5770_ _4137_ _1051_ _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4721_ _4296_ _4299_ _4301_ _4291_ _4302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_124_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7440_ _2577_ _2578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4652_ _4232_ _4233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_30_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7371_ _2417_ _2509_ _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4583_ as2650.cycle\[2\] _4164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5194__I _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9110_ _0003_ clknet_leaf_68_wb_clk_i as2650.r123\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6322_ _0837_ _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9041_ _1595_ _4071_ _4077_ _3742_ _0275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_118_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6253_ _1509_ _1510_ _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6837__A2 _2019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4848__A1 _4428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5896__I0 _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8039__A1 _3151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5204_ _4396_ _0512_ _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6184_ _1234_ _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5135_ _0442_ _0443_ _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7262__A2 _2401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5066_ _0375_ _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_16_wb_clk_i_I clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8211__A1 _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8825_ _3905_ _3906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5576__A2 _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6773__A1 _1949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5968_ _4427_ _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8756_ _1572_ _0566_ _1518_ _3841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_90_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7707_ net34 net33 _2747_ _2839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4919_ _4498_ _4499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7584__I _2340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5899_ _1159_ _1160_ _1176_ _0034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8687_ _1736_ _3769_ _4435_ _3775_ _3776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_139_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7638_ _1634_ _2772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6525__A1 _1757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7569_ _2703_ _2704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8278__A1 _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9308_ _0201_ clknet_leaf_18_wb_clk_i as2650.cycle\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__9320__CLK clknet_leaf_31_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9239_ _0132_ clknet_leaf_39_wb_clk_i as2650.stack\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_55_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8450__A1 _3250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8450__B2 _2513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5264__A1 _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8202__A1 _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5016__A1 _4453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8811__C _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7494__I _2629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8505__A2 _1618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6516__A1 _4383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5319__A2 _4482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8539__B _3633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6059__B _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8441__A1 _2800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5255__A1 _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5255__B2 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8992__A2 _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6940_ _2145_ _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6871_ _2059_ _2061_ _2081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5189__I as2650.r0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5007__A1 _4330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8744__A2 _1764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8610_ _3492_ _3686_ _3331_ _3702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5822_ _1102_ _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6755__A1 as2650.r0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7952__B1 _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5802__I0 _4344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8541_ _3572_ _3624_ _3628_ _3395_ _3635_ _3636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5753_ _1033_ _1034_ _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_72_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4704_ _4284_ _4285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8472_ _1619_ _2540_ _3504_ _3568_ _3569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5684_ as2650.pc\[9\] _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__9343__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7423_ _4390_ _4360_ _2561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4635_ as2650.ins_reg\[4\] as2650.ins_reg\[6\] as2650.ins_reg\[7\] _4216_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7180__A1 _2305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7354_ _2150_ _4393_ _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_25_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_25_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_116_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4566_ _4146_ _4147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6305_ _1515_ _1562_ _1563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7285_ _0654_ _1253_ _1468_ _2423_ _2424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_143_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8168__C _3272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9024_ _1234_ _1233_ _1466_ _4061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_89_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6236_ _4544_ _1453_ _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5494__A1 _4368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6167_ as2650.stack\[4\]\[14\] _1416_ _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_100_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7235__A2 _2363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8432__A1 _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6038__A3 _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5118_ as2650.stack\[2\]\[10\] _0427_ _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6098_ _1367_ _1283_ _1368_ _1370_ _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XTAP_3517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5246__A1 _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5246__B2 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8983__A2 _2449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5049_ _4520_ _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8808_ _0620_ _3588_ _3890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6746__A1 _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8631__C _3420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8739_ _3144_ _1393_ _3824_ _3088_ _3825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_22_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4731__I _4183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7171__A1 _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7171__B2 as2650.stack\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6658__I _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5562__I _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8671__A1 _2477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8806__C _2514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8094__B _4201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5237__A1 _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9216__CLK clknet_leaf_41_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4906__I _4211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5788__A2 _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8726__A2 _3773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6737__A1 _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9366__CLK clknet_leaf_68_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4641__I _4221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8269__B _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8662__A1 _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7070_ _2138_ _2245_ _2251_ _0130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_141_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5476__A1 _4445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6021_ _1294_ _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_6_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8414__A1 _3395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5228__A1 _4494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4816__I _4396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7972_ _3094_ _3096_ _1686_ _2525_ _3097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6976__A1 _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6923_ _2119_ _2130_ _0104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8732__B _2629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6854_ _2063_ _2039_ _2064_ _2065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout49 net50 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_50_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5805_ _1086_ _0341_ _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6785_ _1968_ _1972_ _1998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5647__I as2650.pc\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7940__A3 _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8524_ _3593_ _3618_ _3619_ _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5736_ _0976_ _1022_ _1024_ _0023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5667_ _0962_ _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8455_ as2650.stack\[3\]\[6\] _1920_ _3386_ as2650.stack\[2\]\[6\] _3552_ _3553_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_136_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8350__B1 _3449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7406_ _0910_ _4528_ _2544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4618_ _4198_ _4199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8386_ _0525_ _3485_ _3486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5598_ _0866_ _4466_ _0901_ _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_117_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7337_ _1341_ _2476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8653__A1 _3724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7456__A2 _4512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7268_ _1321_ _2408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5467__A1 _4354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9239__CLK clknet_leaf_39_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6219_ _1095_ _1242_ _4544_ _4199_ _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_63_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9007_ _3230_ _4040_ _4045_ _4046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7199_ _1464_ _2348_ _2349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_63_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8626__C _3598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8956__A2 _2100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_65 io_oeb[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8708__A2 _3769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_76 io_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6941__I _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_87 io_oeb[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6719__A1 _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5557__I _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5942__A2 _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7144__A1 _2265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4902__B1 _4470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8644__A1 _3393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8644__B2 _3598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5458__A1 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7721__B _2852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8947__A2 _2017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4681__A2 _4261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8108__I _3158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7012__I _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8175__A3 _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6186__A2 _1440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6570_ _1779_ _1787_ _1801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_125_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5521_ _4375_ _0610_ _0825_ _4350_ _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8240_ _1696_ _1681_ _3342_ _3343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_117_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5452_ _0757_ _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7686__A2 _2780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6489__A3 _4419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6298__I _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8171_ _2439_ _3186_ _3275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5383_ _0590_ _0689_ _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_7122_ _2282_ _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7438__A2 _2520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7053_ as2650.r123_2\[3\]\[4\] _2239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5930__I as2650.r123_2\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6004_ _0874_ _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8938__A2 _3961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8018__I _2794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9060__A1 _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6949__A1 _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7955_ _1516_ _3080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_70_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8462__B _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6906_ _2108_ _2114_ _2115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_7886_ _2959_ _2990_ _3013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_51_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6837_ as2650.r123_2\[2\]\[2\] _2019_ _2048_ _1980_ _2049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5377__I _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6177__A2 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6768_ _1713_ _1938_ _1981_ _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_7_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5924__A2 _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_40_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_40_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_8507_ _1549_ _2539_ _3603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8688__I _4219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5719_ _0635_ _4416_ _1009_ _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7126__A1 _2215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6699_ _1919_ _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8438_ _2495_ _3530_ _3532_ _3533_ _3089_ _3535_ _3536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__7677__A2 _2809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8874__A1 _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5326__B _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8369_ _1581_ _0496_ _3468_ _3469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_123_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6001__I _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8626__A1 _2926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6936__I _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8929__A2 _3967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9051__A1 _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7601__A2 _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8372__B _3470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7365__A1 _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5287__I _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8314__B1 _3409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7668__A2 _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5679__A1 _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5679__B2 as2650.r123_2\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6340__A2 _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8547__B _3329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8093__A2 _3204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5750__I as2650.r123_2\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5851__A1 _4388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput6 io_in[5] net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_110_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9042__A1 _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6581__I _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7740_ _2867_ _2871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4952_ _4399_ _4532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5197__I net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7671_ _2555_ _2803_ _2804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4883_ _4456_ _4463_ _4464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_75_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6622_ _1778_ _1845_ _1851_ _1806_ _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_127_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6553_ _1747_ _1776_ _1784_ _1760_ _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
X_9341_ _0234_ clknet_leaf_51_wb_clk_i as2650.stack\[6\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5382__A3 _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5504_ as2650.holding_reg\[7\] _0550_ _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7659__A2 _2790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9272_ _0165_ clknet_leaf_12_wb_clk_i as2650.addr_buff\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6484_ as2650.r123\[0\]\[0\] as2650.r123_2\[0\]\[0\] _4146_ _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_134_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8223_ _2408_ _3327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5435_ _0638_ _0664_ _0716_ _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_133_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8608__A1 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8154_ _1329_ _3259_ _3260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5366_ _0672_ _4142_ _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6756__I _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7105_ as2650.r123\[3\]\[5\] _2274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8084__A2 _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8085_ _3164_ _3196_ _3197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5297_ _0597_ _0598_ _0604_ _4389_ _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_59_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8176__C _4200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6095__A1 _4442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7036_ _2191_ _2214_ _2217_ as2650.stack\[4\]\[4\] _2210_ _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_28_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4645__A2 _4225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__9033__A1 _1476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8987_ _3336_ _4010_ _4026_ _4027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7938_ _2824_ _3063_ _3056_ _3064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_128_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7869_ _2385_ _2984_ _2997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8847__A1 _2305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8698__I1 _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8075__A2 _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5570__I _4184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6086__A1 _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5833__A1 _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9024__A1 _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7586__A1 _2720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7497__I _2632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6010__A1 _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8550__A3 _3594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6561__A2 _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8838__A1 _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7510__A1 _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5220_ _0528_ _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_124_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5521__B1 _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5151_ _0444_ _0459_ _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8066__A2 _3175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6077__A1 _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5082_ _4346_ _0358_ _0391_ _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_110_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8910_ _3963_ _3967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__9015__A1 _3136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8369__A3 _3468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8841_ _2300_ _3904_ _3906_ as2650.stack\[6\]\[4\] _3901_ _3918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_53_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4824__I _4285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5588__B1 _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8772_ _0579_ _3856_ _3245_ _3857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5984_ _0814_ _1252_ _1257_ _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7723_ _1497_ _1683_ _2855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4935_ _4389_ _4515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7654_ _2194_ net1 net10 _2187_ _2787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4866_ _4441_ _4446_ _4447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6605_ _0669_ _1723_ _1817_ _1835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_119_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7585_ _2612_ _2720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5655__I as2650.pc\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4797_ _4230_ _4378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9324_ _0217_ clknet_leaf_29_wb_clk_i as2650.pc\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6536_ _1734_ _1752_ _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_88_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9255_ _0148_ clknet_leaf_50_wb_clk_i as2650.stack\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7501__A1 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7870__I as2650.addr_buff\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6467_ _1690_ _1703_ _1705_ _0073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8206_ _1549_ _3309_ _3310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5418_ _0721_ _0723_ _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_45_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9186_ _0079_ clknet_leaf_73_wb_clk_i as2650.r123_2\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6398_ as2650.stack\[3\]\[12\] _1646_ _1650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6486__I _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8137_ _3243_ _3244_ _3245_ _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5349_ _0654_ _0592_ _0655_ _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8068_ _2384_ _3181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5815__A1 _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9006__A1 _4040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7019_ _2216_ _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9006__B2 _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7568__A1 as2650.addr_buff\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5043__A2 _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8650__B _3526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8517__B1 _3596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8296__A2 _3393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6059__A1 _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5806__A1 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4609__A2 as2650.ins_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7271__A3 _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6345__B _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7955__I _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4793__A1 _4368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4720_ _4300_ _4287_ _4301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4651_ _4224_ _4232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7731__A1 _2824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4582_ as2650.cycle\[7\] as2650.cycle\[6\] as2650.cycle\[5\] as2650.cycle\[4\] _4163_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_7370_ _2410_ _2509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6321_ _1278_ _4314_ _1279_ _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_115_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8287__A2 _3386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6252_ _1238_ _1263_ _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_9040_ _1451_ _4075_ _4071_ _4076_ _4077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_116_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5203_ _0463_ _0511_ _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_88_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8039__A2 _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6183_ _1438_ _1439_ _1441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_130_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5134_ as2650.holding_reg\[3\] _0371_ _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9272__CLK clknet_leaf_12_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5065_ _0374_ _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8824_ _2223_ _0626_ _0901_ _3905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8211__A2 _2794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5025__A2 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8755_ _2477_ _0578_ _3839_ _3840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_55_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5967_ _0469_ _1240_ _4432_ _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_40_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7706_ net54 _2838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_40_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4918_ _4439_ _4498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8686_ _4316_ _3772_ _3774_ _3775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5898_ _1124_ _1161_ _1175_ _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_55_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7637_ _2465_ _2771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4849_ _4429_ _4430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7568_ as2650.addr_buff\[7\] _4266_ _2703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_105_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_1_wb_clk_i_I clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7814__B _2943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9307_ _0200_ clknet_leaf_23_wb_clk_i as2650.cycle\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8278__A2 _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6519_ _1734_ _1752_ _1753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_101_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7499_ _2634_ _2635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9238_ _0131_ clknet_leaf_39_wb_clk_i as2650.stack\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9169_ _0062_ clknet_leaf_48_wb_clk_i as2650.stack\[3\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6149__C _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8645__B _3293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6944__I _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5264__A2 _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8202__A2 _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6213__A1 _4255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8269__A2 _3370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7477__B1 _2611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8539__C _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8441__A2 _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6452__A1 _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8729__B1 _3811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6870_ _2059_ _2061_ _2080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5821_ _1067_ _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7685__I _2485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7952__A1 _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7952__B2 _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8540_ _3076_ _3631_ _3634_ _3095_ _3635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_50_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7618__C _2751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5752_ _4200_ _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4703_ as2650.r0\[0\] _4284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8471_ _3345_ _3567_ _3568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5683_ _0963_ _0976_ _0978_ _0016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7422_ _2472_ _2560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4634_ _4181_ _4215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7353_ _2491_ _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4565_ _4145_ _4146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8449__C _3546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6304_ _1518_ _1543_ _1548_ _1561_ _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_144_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7284_ _4427_ _1240_ _4425_ _2423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_89_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9023_ _1359_ _4059_ _4060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6235_ _4550_ _4341_ _0338_ _4417_ _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
Xclkbuf_leaf_65_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_65_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6691__A1 as2650.stack\[1\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6166_ _1012_ _1418_ _1425_ _0052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5117_ _0426_ _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_58_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8432__A2 _3529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6038__A4 _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6097_ _1369_ _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_3507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5048_ _0351_ _0357_ _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_22_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8983__A3 _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8196__A1 _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8807_ _3838_ _1212_ _3888_ _3889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7943__A1 _3065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6746__A2 _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6999_ _1530_ _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8991__I0 _4029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8738_ _2756_ _0476_ _3823_ _3126_ _3824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_41_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9168__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8499__A2 _3594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8669_ _3757_ _3758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5843__I as2650.r123_2\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8671__A2 _4353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8375__B _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8423__A2 _3366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5237__A2 _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7934__A1 _2551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6737__A2 _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4748__A1 _4323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7454__B _2467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5173__A1 _4509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8111__A1 _3164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8662__A2 _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5476__A2 _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6020_ _1293_ _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input4_I io_in[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7971_ net51 _1277_ _3095_ _3096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_66_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6976__A2 _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6922_ _1727_ _2129_ _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4987__A1 _4257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8178__A1 _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9310__CLK clknet_leaf_18_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6853_ _2008_ _2059_ _2064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_62_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7925__A1 _1480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5804_ _4170_ _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6784_ _1968_ _1972_ _1997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8523_ _1391_ _3619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5735_ as2650.stack\[5\]\[8\] _1023_ _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8454_ _3551_ _3552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5666_ _0961_ _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7405_ as2650.pc\[0\] net6 _2543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4617_ _4197_ _4135_ _4198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_50_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8385_ as2650.stack\[4\]\[4\] _3319_ _3322_ as2650.stack\[6\]\[4\] _3320_ as2650.stack\[5\]\[4\]
+ _3485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_50_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5597_ _0900_ _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7336_ _1550_ _2474_ _2475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8102__A1 _3090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7267_ _2406_ _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__8653__A2 _3621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9006_ _4040_ _4034_ _4044_ _1287_ _3230_ _4045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_104_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6218_ _1293_ _0516_ _1229_ _1476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_77_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7198_ _0894_ _2348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8195__B _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6149_ _1397_ _1413_ _1414_ _1410_ _0046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_97_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5219__A2 _4450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4690__A3 _4231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4978__A1 _4348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8169__A1 _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xwrapped_as2650_55 io_oeb[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_66 io_oeb[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_77 io_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xwrapped_as2650_88 io_oeb[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_2669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7916__A1 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4742__I _4160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8341__A1 _3181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5573__I _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8089__C _2624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8884__I _3947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8644__A2 _3727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5458__A2 _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4917__I as2650.r123\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9333__CLK clknet_leaf_80_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7080__A1 _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7907__A1 _2923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4652__I _4232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7168__C _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6186__A3 _1441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5394__A1 _4354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7963__I _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5520_ _4374_ _0824_ _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8332__A1 _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6579__I _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5146__A1 _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5451_ _0756_ _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6343__B1 _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5483__I _4367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6489__A4 _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5697__A2 _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8170_ _3236_ _3273_ _3274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5382_ _0601_ _0599_ _0542_ _0686_ _0688_ _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_7121_ _2280_ _2286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6646__A1 _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7052_ _2238_ _0125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6003_ _1276_ _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5432__B _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8399__A1 _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7203__I _2352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9060__A2 _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6949__A2 _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7954_ _2426_ _3075_ _3078_ _3079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_36_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6905_ _2111_ _2113_ _2114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7885_ as2650.pc\[12\] _0756_ _3012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_78_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4562__I _4142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6836_ _2021_ _2047_ _2048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5385__A1 _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6767_ as2650.r123_2\[2\]\[0\] _1942_ _1979_ _1980_ _1981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7873__I _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8506_ _1709_ _2903_ _3601_ _3602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5718_ _0971_ _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6698_ _1918_ _1919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5137__A1 _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8437_ _4357_ _3345_ _3534_ _3535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__9206__CLK clknet_leaf_73_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5649_ _0946_ _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_80_wb_clk_i clknet_3_0_0_wb_clk_i clknet_leaf_80_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_139_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5688__A2 _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8368_ _3466_ _3439_ _3467_ _3468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_85_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7822__B _2950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7319_ _0717_ _0762_ _2458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XANTENNA__8626__A2 _3706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8299_ _3399_ _3400_ _3401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9356__CLK clknet_leaf_59_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5860__A2 _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9051__A2 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8372__C _3471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7365__A2 _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8562__A1 _3533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8314__A1 _3415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8314__B2 _2549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5679__A2 _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7825__B1 _2952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5300__A1 _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7023__I _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput7 io_in[6] net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XFILLER_49_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9042__A2 _4056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4951_ _4530_ _4531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7670_ _2798_ _2802_ _2803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4882_ as2650.psu\[1\] _4463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8553__A1 _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6621_ _0363_ _1746_ _1763_ _1759_ _1851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_53_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9229__CLK clknet_leaf_62_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7693__I _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9340_ _0233_ clknet_leaf_50_wb_clk_i as2650.stack\[6\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6552_ _4382_ _1748_ _1783_ _4284_ _1784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8305__A1 _2509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5503_ _0544_ _0807_ _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_9271_ _0164_ clknet_leaf_14_wb_clk_i as2650.addr_buff\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6483_ _1718_ _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4590__A2 _4170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6867__A1 _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8222_ _3318_ _3321_ _3325_ _3326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5434_ _0739_ _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__9379__CLK clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8153_ _2484_ _3252_ _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__8608__A2 _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5365_ _0671_ _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6619__A1 _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8457__C _4476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7104_ _2273_ _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8084_ _3194_ _3156_ _3195_ _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5296_ _4397_ _0603_ _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4557__I as2650.ins_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5162__B _4336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6095__A2 _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7292__A1 _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7035_ _2228_ _2229_ _0117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_75_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9033__A2 _4064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7868__I _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8986_ _4012_ _4015_ _4024_ _4025_ _4026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__8792__A1 _3804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7937_ _2686_ _2381_ _3060_ _3062_ _3063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7868_ _2494_ _2996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6819_ _2007_ _2010_ _2031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7799_ _2777_ _2921_ _2929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_74_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8847__A2 _3908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6947__I _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6086__A2 _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7283__A1 _2420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8480__B1 _3576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5294__B1 _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5833__A2 _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9024__A2 _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7586__A2 _2691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8535__A1 _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5349__A1 _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6010__A2 _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4930__I _4509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4572__A2 _4152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8838__A2 _3908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6849__A1 _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7510__A2 _2645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5521__A1 _4375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9380__D _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5521__B2 _4350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5150_ _0413_ _0456_ _0458_ _0407_ _0310_ _0398_ _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai33_1
XFILLER_83_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7274__A1 net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6077__A2 _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5081_ _0383_ _0390_ _4345_ _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_110_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9015__A2 _3216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8840_ _3916_ _3917_ _0234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7577__A2 _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8774__A1 _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5588__A1 _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8771_ _3757_ _3856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5588__B2 _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5983_ _1253_ _1256_ _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7722_ _1479_ _2854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4934_ _4305_ _4306_ _4514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7653_ _2194_ _0682_ _2786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4865_ _4445_ _4446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_127_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4840__I _4190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6604_ _0669_ _1736_ _1817_ _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_14_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7584_ _2340_ _2719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4796_ _4365_ _4376_ _4321_ _4377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_9323_ _0216_ clknet_leaf_24_wb_clk_i as2650.pc\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6535_ _0359_ _1723_ _1751_ _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_105_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5760__A1 _4210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9254_ _0147_ clknet_leaf_50_wb_clk_i as2650.stack\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6466_ _0814_ _1704_ _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4996__B _4310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7501__A2 _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6304__A3 _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8205_ _2754_ _4281_ _3309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5417_ _0640_ _0647_ _0722_ _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_9185_ _0078_ clknet_leaf_73_wb_clk_i as2650.r123_2\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6397_ _1000_ _1643_ _1649_ _0059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8136_ _1565_ _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5348_ _0637_ _0548_ _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7265__A1 _2383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8067_ _3178_ _3179_ _3180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5279_ _0586_ _4141_ _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5815__A2 _4268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7018_ _2215_ _0901_ _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8214__B1 _1638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8765__A1 _3843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8969_ _1570_ _1698_ _4009_ _0271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8517__B2 _3572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7547__B _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6451__B _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5846__I _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4750__I _4257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6677__I _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5503__A1 _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5581__I _4238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7256__A1 net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6059__A2 _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5806__A2 _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7271__A4 _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7008__A1 _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8756__A1 _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6767__B1 _1979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8508__A1 _2334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4650_ _4230_ _4231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput10 io_in[9] net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_128_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4581_ as2650.ins_reg\[3\] _4162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6320_ _1541_ _1536_ _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7192__B _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6251_ _1508_ _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5202_ _0509_ _0510_ _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6182_ _0795_ _0798_ _1438_ _1439_ _1440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_135_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7247__A1 _2383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5133_ as2650.holding_reg\[3\] _0370_ _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_83_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8995__A1 _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8995__B2 _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5064_ _0373_ _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_111_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4835__I _4415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8823_ _3903_ _3904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8754_ _3804_ _0614_ _3839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5966_ _1238_ _1239_ _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7705_ _2830_ _2835_ _2836_ _2837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4917_ as2650.r123\[0\]\[1\] _4497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8685_ _1589_ _3773_ _3774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5981__A1 as2650.psl\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6271__B _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5897_ _1126_ _1174_ _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5666__I _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7636_ _2197_ _2580_ _2769_ _2770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4848_ _4428_ _4136_ _4429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7567_ _2190_ _2686_ _1701_ _2701_ _2702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4779_ _4333_ _4359_ _4360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6930__B1 _2019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9306_ _0199_ clknet_leaf_23_wb_clk_i as2650.cycle\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6518_ _1742_ _1751_ _1752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_106_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7498_ _1532_ _2634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7486__A1 _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9237_ _0130_ clknet_leaf_55_wb_clk_i as2650.stack\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6449_ _1551_ _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_122_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9168_ _0061_ clknet_leaf_48_wb_clk_i as2650.stack\[3\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7238__A1 _4179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8119_ _3208_ _3209_ _3225_ _3228_ _3229_ _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_114_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9099_ _1296_ _3137_ _3135_ _4129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_76_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8986__A1 _4012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7121__I _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8738__A1 _2756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7410__A1 _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6213__A2 _4232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5972__A1 _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6516__A3 _1732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8887__I _3946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7477__A1 _2606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7477__B2 _2613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7229__A1 _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8977__A1 _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5260__B _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6452__A2 _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8729__A1 _3810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8729__B2 _3815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5820_ _1069_ _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7952__A2 _3076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5751_ _4150_ _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5486__I _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4702_ _4282_ _4283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8470_ _1604_ _4370_ _3566_ _3567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_5682_ as2650.stack\[6\]\[8\] _0977_ _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_72_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7421_ _2536_ _2553_ _2554_ _2558_ _2559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4633_ _4162_ _4214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7352_ _1482_ _2481_ _2491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4564_ _4144_ _4145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7468__A1 _2568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6303_ _1547_ _1557_ _1560_ _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_144_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7283_ _2420_ _2421_ _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9022_ _2776_ _1317_ _3282_ _4058_ _4059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__6110__I _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6234_ _1269_ _1237_ _1492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6140__A1 _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8746__B _3831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8417__B1 _3499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6165_ as2650.stack\[4\]\[13\] _1416_ _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_58_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8968__A1 _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5116_ _4459_ _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6096_ _4328_ _1230_ _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5170__B _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7640__A1 _2579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5047_ _0353_ _0355_ _0356_ _0352_ _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_57_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8983__A4 _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8481__B _3577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8806_ _2635_ _0818_ _3887_ _2514_ _3888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6998_ _2193_ _2143_ _2198_ _0111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7943__A2 _3067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8991__I1 _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8737_ _3785_ _0485_ _3822_ _2756_ _3823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5949_ _1089_ _1118_ _4492_ _0792_ _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_55_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8668_ _3746_ _3750_ _3755_ _3756_ _3757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_51_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7619_ _1701_ _2753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5706__A1 _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8599_ _1002_ _3017_ _1599_ _3691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5706__B2 as2650.r123_2\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7459__A1 _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6020__I _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6131__A1 _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6682__A2 _1909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7631__A1 _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6198__A1 _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9112__CLK clknet_leaf_68_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7934__A2 _4187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5945__A1 _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4748__A2 _4328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7698__A1 _2588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9262__CLK clknet_leaf_51_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5173__A2 _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7026__I _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8111__A2 _3221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7970_ _0872_ _3095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6921_ _2122_ _2128_ _2129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_47_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4987__A2 _4386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8178__A2 _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6852_ _2035_ _2038_ _2063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6189__A1 _4311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7925__A2 _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5803_ _4472_ _4484_ _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5397__C1 as2650.stack\[5\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6783_ _1994_ _1995_ _1996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5936__A1 _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8522_ _3210_ _3596_ _3615_ _3617_ _3420_ _3618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5734_ _1021_ _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7689__A1 _2201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8453_ as2650.stack\[0\]\[6\] _3319_ _3320_ as2650.stack\[1\]\[6\] _3551_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__7689__B2 _2681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5665_ _0958_ _0960_ _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7404_ _1336_ _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8350__A2 _3448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4616_ _4196_ _4197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8384_ as2650.stack\[0\]\[4\] _1904_ _1656_ as2650.stack\[1\]\[4\] _3484_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_102_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5596_ _4152_ _0899_ _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_135_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7335_ _2473_ _4361_ _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4911__A2 _4491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8102__A2 _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7266_ _1325_ _2406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6113__A1 _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9005_ _2635_ _3266_ _4041_ _4043_ _4044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7861__A1 _2613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6217_ _1463_ _1467_ _1469_ _1474_ _1475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_132_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7197_ _4393_ _2156_ _2347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4675__A1 _4181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6148_ net21 _1402_ _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_24_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8990__I _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6079_ _1345_ _1351_ _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9135__CLK clknet_leaf_58_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_as2650_56 io_oeb[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8169__A2 _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_67 io_oeb[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_78 io_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_53_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_89 io_oeb[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_96_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7916__A2 _2942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9285__CLK clknet_leaf_27_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6015__I _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8341__A2 _3440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8230__I _3291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8629__B1 _3426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4902__A2 _4482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7852__A1 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4666__A1 _4233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7604__A1 _2588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7080__A2 _2256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5091__A1 as2650.holding_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8405__I _3471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7907__A2 _3029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5918__A1 _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8332__A2 _2641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5450_ _0755_ _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5146__A2 _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6343__A1 as2650.psl\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6343__B2 _4248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_25_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5381_ _4155_ _0687_ _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_2_0_wb_clk_i clknet_0_wb_clk_i clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_7120_ _0912_ _2285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8296__B _3397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8635__A3 _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7843__A1 _2969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7051_ as2650.r123_2\[3\]\[3\] _2238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7843__B2 _2971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9158__CLK clknet_leaf_56_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6002_ _1275_ _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8399__A2 _2762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9060__A3 _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7953_ _1087_ _2441_ _3077_ _3078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_82_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6904_ _2110_ _2112_ _2113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_35_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7884_ _2521_ _3010_ _3011_ _0184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6835_ _2023_ _2046_ _2047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5909__A1 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8571__A2 _3663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_64_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6766_ _1741_ _1980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8505_ _0965_ _1618_ _3601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5717_ as2650.pc\[13\] _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6697_ _4456_ _4458_ _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8323__A2 _3423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8050__I _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5648_ _0945_ _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8436_ _0759_ _2539_ _3534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6334__A1 _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8367_ _0506_ _0366_ _3467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5579_ _4208_ _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7318_ _1316_ _4443_ _0397_ _0339_ _2457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_116_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8298_ _1553_ _4517_ _3400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6098__B1 _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7834__A1 _2895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7249_ _1321_ _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_46_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4648__A1 _4212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4954__S _4333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8653__C _3742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output36_I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5073__A1 _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4753__I _4333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8225__I _3290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4820__A1 _4392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5620__I0 _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7285__B _2423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8314__A2 _3382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8078__A1 _3151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9300__CLK clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5533__B _4231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7825__A1 _2336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9005__B _4041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4639__A1 _4214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput8 io_in[7] net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__7589__B1 _2723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4950_ _4529_ _4530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8002__A1 _4542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4881_ as2650.stack\[2\]\[8\] _4461_ _4462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6620_ _4520_ _1781_ _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5611__I0 _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6551_ _1762_ _1783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5502_ _0794_ _0806_ _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_9270_ _0163_ clknet_leaf_12_wb_clk_i as2650.addr_buff\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6482_ _1716_ _1035_ _1717_ _4202_ _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__6316__A1 _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8221_ as2650.stack\[2\]\[0\] _3322_ _0328_ _3324_ _3325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7923__B _4444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6867__A2 _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5433_ _0636_ _0720_ _0736_ _0738_ _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_127_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5524__C1 _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8738__C _3126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8152_ _1572_ _2477_ _2719_ _3226_ _3258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__8069__A1 _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5364_ as2650.r0\[6\] _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7103_ as2650.r123\[3\]\[4\] _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4838__I _4418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8083_ _2383_ _3061_ _3192_ _3195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7214__I _2357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5295_ _0503_ _0602_ _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_101_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7034_ _0925_ _2224_ _2229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7292__A2 _2408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9033__A3 _4065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8241__A1 _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5055__A1 _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8985_ _3415_ _2438_ _3084_ _3275_ _4025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__8045__I _3157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8792__A2 _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7936_ net26 _1367_ _3061_ _1575_ _1443_ _3062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7867_ _0997_ _2995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_93_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6818_ _2028_ _2029_ _2030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5358__A2 _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7752__B1 _2882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7798_ _2927_ _2928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6749_ _1953_ _1962_ _1963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_137_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9323__CLK clknet_leaf_24_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8419_ as2650.stack\[2\]\[5\] _3518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_87_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7807__A1 _2919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5353__B _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8480__A1 _2526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6086__A3 _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8480__B2 _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5294__B2 _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9024__A3 _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5579__I _4208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8783__A2 _3866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6546__A1 _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5349__A2 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6849__A2 _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7462__C _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5521__A2 _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5809__B1 _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6077__A3 _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8471__A1 _3345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7274__A2 _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5080_ _4354_ _0389_ _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8774__A2 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5982_ _1254_ _1255_ _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_8770_ _3842_ _3854_ _3855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7721_ net54 _2644_ _2852_ _2853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4933_ _4511_ _4512_ _4513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_75_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7652_ _2636_ _2760_ _2696_ _2726_ _2785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_4864_ _4415_ _4444_ _4445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9346__CLK clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6603_ _1830_ _1831_ _1832_ _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7583_ _2695_ _2717_ _2718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_53_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4795_ _4375_ _4376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7209__I _2357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_59_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_59_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_9322_ _0215_ clknet_leaf_29_wb_clk_i as2650.pc\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6534_ _1756_ _1766_ _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_53_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5760__A2 _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8749__B _3757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9253_ _0146_ clknet_leaf_55_wb_clk_i as2650.stack\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6465_ _1697_ _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6304__A4 _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8204_ _3093_ _3300_ _3307_ _3308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5416_ _0659_ _0653_ _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9184_ _0077_ clknet_leaf_69_wb_clk_i as2650.r123_2\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6396_ as2650.stack\[3\]\[11\] _1646_ _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_47_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8135_ _1486_ _0893_ _3209_ _1507_ _3244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__4568__I _4148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5347_ _0414_ _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_47_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8066_ _0687_ _3175_ _3179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8462__A1 _2201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7265__A2 _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5278_ _0585_ _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7017_ _4474_ _2215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5815__A3 _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8214__A1 as2650.stack\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8765__A2 _3848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8968_ _2373_ _1704_ _4009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7828__B _2661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7919_ _1320_ _3045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8899_ _1674_ _3949_ _3957_ _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5200__A1 _4218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8659__B _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6958__I _2163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7789__I net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5267__A1 _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9219__CLK clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8205__A1 _2754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7008__A2 _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5019__A1 as2650.stack\[7\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8756__A2 _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9369__CLK clknet_leaf_74_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6767__B2 _1980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8508__A2 _2755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4941__I _4286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7192__A1 _2150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4580_ _4157_ _4160_ _4161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5742__A2 _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8569__B _3662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5772__I _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6250_ _1346_ _1507_ _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_115_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8692__A1 _3767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5201_ _4533_ _4524_ _4510_ _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6181_ as2650.psl\[1\] _0795_ _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7247__A2 _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5132_ as2650.r123\[0\]\[3\] _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5063_ net8 _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8747__A2 _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8822_ _0958_ _2212_ _3903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_4_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8753_ _2386_ _3838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5965_ _4136_ _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_40_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7704_ _1330_ _2836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4916_ _4275_ _4414_ _4496_ _0000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5896_ _0570_ _1173_ _1145_ _1174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_55_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8684_ _3771_ _3773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5981__A2 _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7635_ _2752_ _2768_ _2573_ _2769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4847_ _4197_ _4428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_7566_ _2693_ _2700_ _1252_ _2701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4778_ _4356_ _4358_ _4359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6930__A1 _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9305_ _0198_ clknet_3_3_0_wb_clk_i as2650.halted vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_140_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6517_ _1743_ _1747_ _1750_ _1751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_140_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7497_ _2632_ _2633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9236_ _0129_ clknet_leaf_64_wb_clk_i as2650.r123_2\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6448_ _1689_ _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9167_ _0060_ clknet_leaf_49_wb_clk_i as2650.stack\[3\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6379_ _1611_ _1515_ _1635_ _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8118_ _1301_ _3229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6727__B _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9098_ as2650.psu\[4\] _4127_ _4128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5249__B2 _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8986__A2 _4015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8049_ _1354_ _2348_ _3162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7402__I _2539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6997__A1 _2197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5350__C _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8738__A2 _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6018__I _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7558__B _2502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8233__I _2387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5972__A2 _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7174__A1 _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6516__A4 _1749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4932__B1 _4507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5592__I _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7229__A2 _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4936__I _4147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8977__A2 _3773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9191__CLK clknet_leaf_47_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8729__A2 _4388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7937__B1 _3060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6372__B _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__9386__D _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8143__I _4171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5750_ as2650.r123_2\[0\]\[0\] _1032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_76_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4701_ _4280_ _4281_ _4282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5681_ _0962_ _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7982__I _1486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7420_ _2555_ _2557_ _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4632_ _4195_ _4212_ _4213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5715__A2 _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7351_ _1311_ _2478_ _2489_ _2490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4563_ as2650.psl\[4\] _4144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_128_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6302_ _1558_ _1291_ _1559_ _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_144_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8665__A1 _1939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7282_ _4551_ _1501_ _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5479__A1 _4274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6233_ _1490_ _1317_ _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9021_ _4491_ _3268_ _2404_ _4057_ _4058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__6140__A2 _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8746__C _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8417__A1 _3250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6164_ _1006_ _1418_ _1424_ _0051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8417__B2 _2513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5115_ as2650.stack\[3\]\[10\] _4452_ _4454_ _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8968__A2 _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8318__I _3376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9090__A1 _4065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6095_ _4442_ _1228_ _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__7222__I _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5046_ _0349_ _4505_ _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_38_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8481__C _3076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8196__A3 _3299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8805_ _3785_ _0828_ _3182_ _3886_ _3887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_53_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5677__I _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6997_ _2197_ _2164_ _2168_ as2650.stack\[2\]\[5\] _2142_ _2198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
Xclkbuf_leaf_74_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_74_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4581__I as2650.ins_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8736_ _2338_ _0491_ _3822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_40_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5948_ _1212_ _1083_ _1222_ _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_107_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8667_ _1318_ _1476_ _1478_ _1484_ _3756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_139_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5879_ _1124_ _1144_ _1157_ _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_55_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7618_ _2719_ _2731_ _2750_ _2751_ _2752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_107_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6903__A1 _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8598_ _3394_ _3688_ _3689_ _3471_ _3690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7549_ _2517_ _2684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6301__I _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7459__A2 _2592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8656__A1 _2755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8656__B2 _3175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9219_ _0112_ clknet_leaf_54_wb_clk_i as2650.stack\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6131__A2 _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8656__C _4260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5890__A1 _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9081__A1 _4113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8672__B _3080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5642__A1 as2650.stack\[5\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7934__A3 _3059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5945__A2 _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7147__A1 _2305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8344__B1 _3433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7147__B2 as2650.stack\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7698__A2 _2828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8895__A1 _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_15_wb_clk_i_I clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9008__B _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8647__A1 _3724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5255__C _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6122__A2 _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9072__A1 _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8582__B _3441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6920_ _2123_ _2127_ _2128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_130_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6851_ _2059_ _2060_ _2061_ _2062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_1_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6189__A2 _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5802_ _4344_ _1081_ _1083_ _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5397__B1 _4466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_54_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5397__C2 _4470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6782_ _1992_ _1993_ _1995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8521_ _1085_ _1499_ _3046_ _3616_ _3617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5733_ _1021_ _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7689__A2 _2684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8452_ _0947_ _3529_ _3550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_104_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8886__A1 _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5664_ _0959_ _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7403_ _2530_ _2532_ _2535_ _2536_ _2537_ _2540_ _2541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_135_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4615_ _4138_ _4196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5595_ _0873_ _0875_ _0892_ _0897_ _0898_ _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_8383_ as2650.stack\[2\]\[4\] _1639_ _3483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6121__I _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7334_ _2472_ _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8638__A1 _4264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5165__C _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7265_ _2383_ _1547_ _2404_ _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_46_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7310__A1 _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5960__I _4443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9004_ _4042_ _4030_ _1009_ _3123_ _0619_ _4043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__5321__B1 _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6216_ _1045_ _1470_ _1473_ _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__7861__A2 _2984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7196_ _1500_ _1349_ _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_63_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5872__A1 _4527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4675__A2 _4255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9063__A1 _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6147_ _1411_ _1398_ _1412_ _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7613__A2 _2690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6078_ _1347_ _1350_ _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8810__A1 _3262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5029_ _4277_ _4423_ _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_73_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4978__A3 _4506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_as2650_57 io_oeb[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8169__A3 _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_68 io_oeb[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_96_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xwrapped_as2650_79 io_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__7377__A1 _2490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8719_ _3804_ _2592_ _3805_ _3806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7129__A1 _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8877__A1 _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8629__A1 _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8629__B2 _3706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6966__I _2163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7301__A1 _4431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7852__A2 _2942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4666__A2 _4206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9054__A1 _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7604__A2 _2735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8801__A1 _2458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7797__I _2855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4969__A3 _4548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5091__A2 _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6206__I _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6040__A1 _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7540__A1 _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6343__A2 _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5380_ _4182_ _4193_ _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_126_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8635__A4 _3663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7050_ _2237_ _0124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5713__C _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7843__A2 _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6001_ _0879_ _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_95_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__9060__A4 _2631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7952_ _2396_ _3076_ _2407_ _1163_ _1319_ _3077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_54_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5082__A2 _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6903_ _0788_ _2084_ _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7883_ _2982_ _2942_ _2943_ _3011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7359__A1 _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6834_ _1994_ _2045_ _2046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_62_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5909__A2 _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6765_ _1944_ _1978_ _1979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_50_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6582__A2 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5955__I _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8504_ _3103_ _3598_ _3353_ _3599_ _3600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_5716_ _0977_ _1006_ _1007_ _0020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_91_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6696_ _1674_ _1909_ _1917_ _0090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8435_ _2645_ _3533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5647_ as2650.pc\[6\] _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7531__A1 _2584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6334__A2 _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8366_ _0506_ _0366_ _3466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5578_ _4254_ _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7317_ _2428_ _2430_ _2431_ _2455_ _2456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__5690__I _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8297_ _0373_ _4517_ _3399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6098__A1 _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6098__B2 _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7248_ _1367_ _1279_ _2346_ _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8492__C1 _3588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5845__A1 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4648__A2 _4228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9036__A1 _4072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7179_ _2199_ _2311_ _2330_ _0160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_58_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7598__A1 _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9252__CLK clknet_leaf_63_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6270__A1 _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6022__A1 _4199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7566__B _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7770__A1 _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5620__I1 as2650.stack\[5\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4584__A1 as2650.cycle\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4887__A2 _4458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8078__A2 _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6089__A1 _4394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7825__A2 _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9005__C _4043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4639__A2 _4219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9027__A1 _1475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7038__B1 _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7589__A1 _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput9 io_in[8] net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XANTENNA__7589__B2 _2681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8002__A2 _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4880_ _4460_ _4461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5775__I _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7761__A1 _2788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5611__I1 as2650.stack\[5\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8151__I _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6550_ _4285_ _1781_ _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_140_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5501_ _0719_ _0727_ _0805_ _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6481_ _1714_ _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__6316__A2 _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8220_ _3323_ _3324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5432_ _0565_ _0737_ _0636_ _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_127_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4878__A2 _4458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8151_ _3256_ _3257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8069__A2 _3181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5363_ _0669_ _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8100__B _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7102_ _2272_ _0141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8082_ _1685_ _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5294_ _0509_ _0463_ _0599_ _0601_ _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_141_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5827__A1 _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7033_ _2183_ _2219_ _2220_ as2650.stack\[4\]\[3\] _2221_ _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_113_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5015__I _4478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8777__B1 _3184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4854__I _4434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8241__A2 _3181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8984_ _1046_ _4020_ _4022_ _4023_ _4024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6252__A1 _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7935_ _1324_ _3061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7866_ _2719_ _2993_ _2483_ _2994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_93_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6817_ _0750_ _2027_ _2002_ _2029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_23_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7752__A1 _2467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7797_ _2855_ _2927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6555__A2 _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5685__I _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7752__B2 _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6748_ as2650.r0\[6\] _1744_ _1962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6679_ _1906_ _1907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8418_ _3515_ _3516_ _3517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9106__B _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8349_ as2650.stack\[7\]\[3\] _1919_ _1638_ as2650.stack\[6\]\[3\] _4475_ _3450_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_133_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7807__A2 _2644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8480__A2 _3562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8768__B1 _3850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4764__I _4247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6243__A1 _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5046__A2 _4505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7991__A1 _4406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6546__A2 _1749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9148__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4939__I as2650.r0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5809__A1 _4295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6482__A1 _1716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4674__I as2650.ins_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5981_ as2650.psl\[7\] _1239_ _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_65_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7720_ _1516_ _2851_ _2852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4932_ _4502_ _4504_ _4507_ _4510_ _4512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__4796__A1 _4365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7651_ _2783_ _2784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_75_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4863_ _4443_ _4426_ _4444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__7734__A1 _2774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6602_ _1801_ _1820_ _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_21_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7582_ _2636_ _2659_ _2716_ _2717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4794_ _4374_ _4375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9321_ _0214_ clknet_leaf_31_wb_clk_i as2650.pc\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6533_ _1758_ _1760_ _1765_ _1766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_118_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8749__C _3834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9252_ _0145_ clknet_leaf_63_wb_clk_i as2650.r123\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6464_ _1292_ _1692_ _1702_ _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8203_ _4161_ _3304_ _3306_ _1251_ _3307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5415_ _0719_ _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_9183_ _0076_ clknet_leaf_74_wb_clk_i as2650.r123_2\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6395_ _0993_ _1643_ _1648_ _0058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_leaf_28_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_28_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_82_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8134_ as2650.cycle\[4\] _3243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5346_ _4421_ _0591_ _0652_ _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_82_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8065_ _1342_ _3178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8462__A2 _3377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5277_ as2650.r0\[5\] _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5276__A2 _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7016_ _2213_ _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8214__A2 _1919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6225__A1 _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8967_ _3191_ _1698_ _4008_ _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_37_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4787__A1 _4367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7918_ _2445_ _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_93_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8898_ as2650.stack\[7\]\[14\] _3947_ _3957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_62_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7849_ net53 _1711_ _2851_ _2977_ _2978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_51_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7725__A1 _2648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5200__A2 _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7135__I _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4711__A1 _4291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8438__C1 _3089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8453__A2 _3319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8394__C _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6464__A1 _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5267__A2 _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8205__A2 _4281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6216__A1 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6767__A2 _1942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7192__A2 _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8569__C _3592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8141__A1 _2416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4669__I _4249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8692__A2 _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5200_ _4218_ _0355_ _4507_ _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_131_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6180_ _0810_ _1431_ _1437_ _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5131_ _0347_ _4499_ _0440_ _0002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_83_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7247__A3 _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5062_ _0371_ _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6207__A1 _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9313__CLK clknet_leaf_18_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8821_ _3901_ _3902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8752_ _3763_ _3837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5964_ _4197_ _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7703_ _2704_ _2833_ _2834_ _2476_ _2835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_40_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4915_ as2650.r123\[0\]\[0\] _4440_ _4495_ _4496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8683_ _3771_ _3772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7707__A1 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5895_ _0614_ _1060_ _1172_ _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7634_ _2196_ _2686_ _2753_ _2767_ _2768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4846_ _4421_ _4427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8380__A1 _3458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8380__B2 _3291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7565_ _2687_ _1710_ _2500_ _2699_ _2700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_105_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4777_ _4357_ as2650.addr_buff\[5\] _4358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5963__I _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6930__A2 _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9304_ _0197_ clknet_3_0_0_wb_clk_i as2650.holding_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6516_ _4383_ _4294_ _1732_ _1749_ _1750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_14_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8132__A1 _2633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7496_ _2631_ _2632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9235_ _0128_ clknet_leaf_62_wb_clk_i as2650.r123_2\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4579__I _4159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6447_ _1688_ _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6694__A1 _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9166_ _0059_ clknet_leaf_48_wb_clk_i as2650.stack\[3\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6378_ _1634_ _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_103_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8117_ _3226_ _3227_ _3207_ _3228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_62_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5329_ _0395_ _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_62_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9097_ _2373_ _3144_ _4121_ _4127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6446__A1 _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6727__C _4438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8048_ _3156_ _3160_ _3059_ _3161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_130_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8199__A1 _2458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7946__A1 _4237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8371__A1 _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5724__A3 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8123__A1 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4932__B2 _4510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4791__S0 _4197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8426__A2 _3524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9080__I _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9336__CLK clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7634__B1 _2753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4999__A1 _4302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7937__A1 _2686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4952__I _4399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_44_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4700_ as2650.r123\[2\]\[0\] as2650.r123_2\[2\]\[0\] _4147_ _4281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5680_ _0975_ _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7165__A2 _2248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4631_ _4206_ _4211_ _4212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7350_ _2418_ _2480_ _2483_ _2488_ _2489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_15_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4562_ _4142_ _4143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8114__A1 _3210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6301_ _1526_ _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8665__A2 _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7281_ _0654_ _1493_ _2419_ _2420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_143_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5479__A2 _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9020_ _0553_ _1364_ _4057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6232_ _1489_ _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8417__A2 _3495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6163_ as2650.stack\[4\]\[12\] _1420_ _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5114_ _4276_ _0392_ _0423_ _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6094_ _4194_ _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6119__I _4202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5045_ _0354_ _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_22_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7928__A1 _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4862__I _4442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8804_ _2338_ _0830_ _3886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6996_ _2196_ _2197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5403__A2 _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8735_ _3703_ _3821_ _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5947_ _1083_ _1221_ _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8666_ _1333_ _1474_ _3753_ _3754_ _3755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__8353__A1 _3333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5878_ _1126_ _1156_ _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7156__A2 _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7617_ _2483_ _2751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4829_ _4363_ _4404_ _4409_ _4410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8597_ _3020_ _3669_ _3689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6903__A2 _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7548_ _2579_ _2682_ _2683_ _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7479_ _2540_ _2611_ _2616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8656__A2 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9359__CLK clknet_leaf_59_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9218_ _0111_ clknet_leaf_56_wb_clk_i as2650.stack\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9149_ _0042_ clknet_leaf_15_wb_clk_i net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8408__A2 _3468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7413__I _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7616__B1 _2749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5890__A2 _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9081__A2 _4100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7092__A1 _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7092__B2 as2650.stack\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5642__A2 _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5868__I _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4772__I _4352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8592__A1 as2650.pc\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8344__A1 _3415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7147__A2 _2286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8344__B2 _2524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6699__I _1919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8895__A2 _3949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4721__B _4291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4905__A1 _4472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8647__A2 _3148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5108__I _4330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8847__C _3900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4947__I _4526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9072__A2 _3144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7083__A1 _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6830__A1 _2001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5778__I _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6850_ _0585_ _1970_ _2061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8583__A1 _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5801_ _1082_ _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5397__A1 as2650.stack\[7\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6781_ _1992_ _1993_ _1994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5397__B2 as2650.stack\[4\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8520_ _3426_ _3596_ _3616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5732_ _1020_ _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8335__A1 _2793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8451_ _3153_ _3547_ _3548_ _3549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5149__A1 _4518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5663_ _0856_ _0900_ _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8886__A2 _3948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7402_ _2539_ _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4614_ _4191_ _4194_ _4195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_102_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8382_ as2650.stack\[3\]\[4\] _2215_ _4473_ _3482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_141_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5594_ _0891_ _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7333_ _4267_ _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8638__A2 _3158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5018__I _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7264_ _1282_ _1361_ _2404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7310__A2 _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9003_ _1921_ _1640_ _4042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4857__I _4202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6215_ _1471_ _0394_ _1472_ _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_89_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7195_ _1086_ _1683_ _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_131_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6146_ _1399_ _0754_ _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9063__A2 _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7074__A1 _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7074__B2 as2650.stack\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6077_ _0883_ _1315_ _1349_ _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_100_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8810__A2 _3793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5028_ _0338_ _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA_input10_I io_in[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4592__I as2650.cycle\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4978__A4 _4509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8169__A4 _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_58 io_oeb[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_69 io_oeb[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_54_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7377__A2 _2515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5388__A1 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6979_ _2181_ _2182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8718_ _3785_ _0358_ _3805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8326__A1 _2181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7129__A2 _2286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8649_ _0781_ _3327_ _2388_ _3727_ _3739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_142_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6312__I _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6888__A1 _2021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4899__B1 _4461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7852__B _2943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8629__A2 _3481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7301__A2 _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4666__A3 _4242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9054__A2 _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8262__B1 _3362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8801__A2 _2753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8565__A1 _3250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8565__B2 _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6040__A2 _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8702__I _4227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8317__A1 _3329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5551__A1 _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6000_ _1272_ _1273_ _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_80_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input2_I io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5067__B1 _4510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7951_ _2157_ _3076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6902_ _2061_ _2110_ _2086_ _2087_ _2111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_78_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7882_ _0997_ _2522_ _3009_ _2940_ _3010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_39_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8556__A1 _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7359__A2 _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6833_ _2026_ _2044_ _2045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_51_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8612__I _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6764_ _1947_ _1977_ _1978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_11_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8308__A1 _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8503_ _2204_ _3570_ _0965_ _3599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5715_ as2650.stack\[6\]\[12\] _0986_ _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6695_ as2650.stack\[1\]\[14\] _1907_ _1917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_13_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8434_ _1709_ _2790_ _3531_ _3532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5646_ _0752_ _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7531__A2 _2585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7672__B _2467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8365_ _3256_ _3457_ _3464_ _2524_ _2927_ _3465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5577_ as2650.addr_buff\[7\] _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8487__C _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7316_ _2445_ _2447_ _2454_ _2455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_8296_ _3382_ _3393_ _3397_ _3398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6098__A2 _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4587__I as2650.cycle\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7295__A1 _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7247_ _2383_ _2386_ _2380_ _2388_ _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_137_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8492__C2 _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7178_ _2265_ _2313_ _2316_ as2650.stack\[0\]\[6\] _2320_ _2330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__9036__A2 _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6129_ _1375_ _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5058__B1 _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7598__A2 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6270__A2 _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6022__A2 _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7770__A2 _2886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7138__I _2190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6042__I _4232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5533__A1 _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5881__I as2650.r123_2\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6198__B _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7286__A1 _2419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6089__A2 _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7038__A1 _2197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7589__A2 _2684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8786__A1 _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8538__A1 _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7210__A1 _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5221__B1 _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5500_ _0737_ _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6480_ _0853_ _4489_ _1716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8710__A1 _3791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5431_ _0730_ _0718_ _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5524__A1 _4375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5524__B2 _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8150_ _2437_ _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5362_ _0586_ _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7101_ as2650.r123\[3\]\[3\] _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8081_ _3191_ _3192_ _3067_ _3154_ _3193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_142_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5293_ _4155_ _0600_ _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7032_ _2226_ _2227_ _0116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_141_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8777__A1 _3838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8983_ _3844_ _2449_ _1281_ _1357_ _4023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_83_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7934_ _2551_ _4187_ _3059_ _3060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_43_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5031__I _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7865_ _2990_ _2992_ _2993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_36_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7201__A1 _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6816_ _2027_ _2002_ _2028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7796_ _2925_ _2926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7752__A2 _2874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6747_ as2650.r0\[7\] _1730_ _1961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5763__A1 _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6678_ _0866_ _1905_ _0960_ _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__8701__A1 _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8417_ _3250_ _3495_ _3499_ _2513_ _3154_ _3516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__5515__A1 _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5629_ _0928_ _0903_ _0929_ _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8348_ as2650.stack\[4\]\[3\] _1903_ _1655_ as2650.stack\[5\]\[3\] _3449_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_117_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8279_ _0919_ _3380_ _3381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_132_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8768__A1 _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8768__B2 _3852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6243__A2 _4167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7991__A2 _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5754__A1 _4248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5506__A1 _4336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7259__A1 _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8456__B1 _3386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5809__A2 _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6482__A2 _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8427__I _3290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7431__A1 _2568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6234__A2 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5980_ as2650.psl\[6\] _4428_ _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_92_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8590__C _3331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4931_ _4502_ _4504_ _4507_ _4510_ _4511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XTAP_3490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5993__A1 _4174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4796__A2 _4376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5786__I _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7650_ as2650.pc\[6\] net2 _2783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_127_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4862_ _4442_ _4443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6601_ _1801_ _1820_ _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_20_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7581_ _2181_ _0507_ _2716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5745__A1 _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4793_ _4368_ _4371_ _4373_ _4374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_9320_ _0213_ clknet_leaf_31_wb_clk_i as2650.pc\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6532_ _4405_ _1764_ _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9251_ _0144_ clknet_leaf_63_wb_clk_i as2650.r123\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6463_ _1502_ _1701_ _1702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9242__CLK clknet_leaf_55_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8111__B _3067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8202_ _0864_ _2440_ _3305_ _4161_ _3306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_118_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6410__I _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5414_ _0719_ _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6170__A1 _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9182_ _0075_ clknet_leaf_8_wb_clk_i as2650.ins_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6394_ as2650.stack\[3\]\[10\] _1646_ _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8133_ _3151_ _0893_ _3235_ _3242_ _3229_ _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_115_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5345_ as2650.holding_reg\[5\] _4191_ _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4720__A2 _4287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5026__I _4542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8765__C _3767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8998__A1 _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8064_ _1354_ _3175_ _2390_ _3176_ _3177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5276_ _4298_ _0583_ _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_68_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_68_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4865__I _4445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7015_ _0622_ _2212_ _2213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_130_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7241__I _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8966_ _1556_ _1704_ _4008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7973__A2 _3097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7917_ _2521_ _3042_ _3043_ _0185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_110_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5696__I _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4787__A2 _4142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5984__A1 _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8897_ _1672_ _3949_ _3956_ _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_93_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7848_ _1546_ _2976_ _2977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5736__A1 _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7779_ _2884_ _2771_ _2772_ _2910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5200__A3 _4507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7844__C _2551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7489__A1 _2615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7416__I _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8438__C2 _3535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4711__A2 _4190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8989__A1 _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6464__A2 _1692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6216__A2 _1470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9115__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5539__C _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8913__A1 _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5727__A1 as2650.stack\[6\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9265__CLK clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7326__I _2464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8585__C _2927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5130_ _4500_ _0424_ _0439_ _4498_ _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_97_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7247__A4 _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7652__A1 _2636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_73_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8157__I as2650.psu\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5061_ _0370_ _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6207__A2 _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8820_ _3900_ _3901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5966__A1 _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8751_ _3189_ _3836_ _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5963_ _0854_ _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_80_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7702_ _1680_ _2704_ _2834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4914_ _4439_ _4447_ _4486_ _4494_ _4495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_5894_ _1136_ _1170_ _1171_ _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_8682_ _0550_ _3770_ _0340_ _3771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__7707__A2 net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7633_ _0940_ _2655_ _2766_ _1443_ _2767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_21_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4845_ _4420_ _4422_ _4425_ _4426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_138_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8380__A2 _3457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7564_ _1545_ _2698_ _2699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4776_ as2650.addr_buff\[6\] _4357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_119_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6515_ _1748_ _1749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9303_ _0196_ clknet_leaf_2_wb_clk_i as2650.holding_reg\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_119_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7495_ _2443_ _2631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8132__A2 _3237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6446_ _1677_ _1118_ _1356_ _1687_ _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
X_9234_ _0127_ clknet_leaf_62_wb_clk_i as2650.r123_2\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8776__B _2514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7680__B _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7891__A1 _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6694__A2 _1909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9165_ _0058_ clknet_leaf_48_wb_clk_i as2650.stack\[3\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6377_ _1565_ _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8116_ _1429_ _1493_ _1494_ _3220_ _3227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_5328_ as2650.r123\[0\]\[5\] _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9096_ _4122_ _4124_ _4126_ _3249_ _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_138_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6446__A2 _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8047_ _3158_ _3159_ _3160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5259_ as2650.holding_reg\[4\] _0566_ _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8986__A4 _4025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9138__CLK clknet_leaf_46_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8199__A2 _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7946__A2 _2348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9288__CLK clknet_leaf_27_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8949_ _0424_ _3992_ _3993_ as2650.r123\[2\]\[2\] _3997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5957__A1 _4219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6315__I _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5709__A1 _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8371__A2 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7146__I _2204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6050__I _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7590__B _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7882__A1 _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7882__B2 _2940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4791__S1 _4148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7634__A1 _2196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8831__B1 _3909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8705__I _3792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7937__A2 _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5948__A1 _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7765__B _2607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4630_ _4210_ _4211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_50_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6373__A1 _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6373__B2 _1627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4561_ _4141_ _4142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6300_ _0597_ _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7280_ _4199_ _4544_ _2419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6125__A1 _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8665__A3 _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6231_ _0882_ _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4687__A1 _4263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6162_ _1000_ _1417_ _1423_ _0050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_135_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7625__A1 _2756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5113_ _4276_ _0422_ _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6093_ _1359_ _1365_ _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5044_ _0349_ _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5100__A2 _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8615__I _3705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7928__A2 _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8803_ _3837_ _3884_ _3885_ _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5939__A1 _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6995_ _2195_ _2196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8734_ _0917_ _3758_ _3820_ _3821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5946_ _0828_ _1057_ _1220_ _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8665_ _1939_ _0871_ _1352_ _1487_ _3754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_5877_ _1145_ _1154_ _1155_ _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__8353__A2 _3425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7616_ _2661_ _2746_ _2749_ _2480_ _2658_ _2750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4828_ _4406_ _4362_ _4408_ _4409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6364__A1 _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8596_ _1003_ _3687_ _3688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6364__B2 _1611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7547_ _2643_ _2466_ _1635_ _2683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4759_ _4319_ _4327_ _4339_ _4340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_135_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7478_ _1337_ _2600_ _2614_ _2615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5923__B _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9217_ _0110_ clknet_leaf_53_wb_clk_i as2650.stack\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6429_ as2650.stack\[2\]\[13\] _1659_ _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_136_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4678__A1 _4198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_12_wb_clk_i clknet_3_2_0_wb_clk_i clknet_leaf_12_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5875__B1 _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9148_ _0041_ clknet_leaf_15_wb_clk_i net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7616__A1 _2661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7616__B2 _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9079_ _4365_ _4111_ _4112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8592__A2 _3663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8344__A2 _3424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4905__A2 _4484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9091__I _4121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7083__A2 _2256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5094__A1 _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8435__I _2645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8583__A2 _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5800_ _1047_ _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6780_ _0586_ _1887_ _1993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5731_ _1018_ _1019_ _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_95_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8450_ _3250_ _3530_ _3532_ _2513_ _3154_ _3548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_31_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5149__A2 _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5662_ _0957_ _0430_ _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6346__A1 _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7401_ _2538_ _2539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4613_ _4156_ _4192_ _4193_ _4194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_8381_ _2391_ _3481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5593_ _0447_ _0896_ _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7332_ _1550_ _2470_ _2471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_128_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7846__A1 _2961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7263_ _1327_ _2403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6214_ _4433_ _4489_ _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7310__A3 _4425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9002_ _3122_ _4041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7194_ _1351_ _2341_ _2342_ _2343_ _2344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__5321__A2 _4482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6145_ _0790_ _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6076_ as2650.cycle\[3\] _1348_ _4174_ _4172_ _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5085__A1 _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4873__I _4453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5027_ _4420_ _4488_ _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8023__A1 _2736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_59 io_oeb[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6585__A1 _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5388__A2 _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6978_ as2650.pc\[3\] _2181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6585__B2 _1757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8717_ _2337_ _3804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5929_ _1192_ _1160_ _1204_ _0036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8326__A2 _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9326__CLK clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8648_ _3214_ _3735_ _3737_ _3738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8579_ _3459_ _3667_ _3670_ _3504_ _3671_ _3672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_108_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7837__A1 _2658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8964__B _3962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4666__A4 _4246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8262__B2 as2650.stack\[5\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5076__A1 _4357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4783__I _4221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8014__A1 _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6576__A1 _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5379__A2 _4506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8317__A2 _3382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5119__I _4465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5000__A1 _4302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5551__A2 _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4958__I _4221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7334__I _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8253__A1 _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5067__A1 _4218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5067__B2 _4533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7950_ _2450_ _3074_ _2412_ _2451_ _3075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6901_ _0750_ _2109_ _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7002__C _2173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7881_ _2989_ _2994_ _3003_ _3008_ _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_78_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8556__A2 _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6832_ _2030_ _2043_ _2044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_62_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9349__CLK clknet_leaf_51_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6763_ _1949_ _1976_ _1977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_50_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7509__I _2352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8308__A2 _2754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8502_ _3057_ _3598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5714_ _1005_ _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7516__B1 _2651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6694_ _1672_ _1909_ _1916_ _0089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8433_ _0946_ _1618_ _3531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5645_ _0938_ _0861_ _0943_ _0013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8768__C _1513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7672__C _2804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8364_ _1679_ _2698_ _3463_ _3464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5576_ _0877_ _0879_ _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5542__A2 _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7819__A1 _2744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7315_ _1501_ _1504_ _2351_ _2453_ _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_144_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7244__I _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8295_ _3395_ _3396_ _3397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8492__A1 _3317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7295__A2 _2433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7246_ _2387_ _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7177_ _0938_ _2311_ _2329_ _0159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_131_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6128_ _1372_ _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8244__A1 _3089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5699__I _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5058__B2 _4521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6059_ _1323_ _1324_ _1331_ _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_2_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4805__A1 _4381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6558__A1 _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6323__I _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5533__A2 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8483__A1 _3293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7286__A2 _2424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5297__A1 _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9027__A3 _4060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8235__A1 _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5830__C _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8786__A2 _3766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6549__A1 _4147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5221__A1 as2650.stack\[0\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5221__B2 as2650.stack\[2\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7773__B _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4980__B1 _4506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5430_ _0726_ _0729_ _0735_ _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8710__A2 _3796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5524__A2 _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6721__A1 _4195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5361_ _0667_ _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_103_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7100_ _2271_ _0140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8474__A1 _2203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8080_ _2432_ _3192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5292_ _4182_ _4158_ _4177_ _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_113_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7031_ _0918_ _2224_ _2227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8226__A1 _3316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8777__A2 _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6408__I _1656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8982_ _1498_ _3236_ _4021_ _4022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__9171__CLK clknet_leaf_60_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout53_I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7933_ _3058_ _3059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7864_ _2991_ _2965_ _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6815_ _1887_ _2027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5212__A1 _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7795_ _1479_ _2925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6143__I _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6746_ _1879_ _1885_ _1959_ _1960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4799__S _4379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6677_ _1904_ _1905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8701__A2 _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8416_ _3497_ _3514_ _3391_ _3515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6712__A1 as2650.stack\[0\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5628_ as2650.stack\[5\]\[3\] _0904_ _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8347_ as2650.stack\[0\]\[3\] _1903_ _1655_ as2650.stack\[1\]\[3\] _0328_ _3448_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5559_ _0862_ _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_133_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8465__A1 _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8278_ _0910_ _0862_ _3380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5279__A1 _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5931__B _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7229_ _2372_ _2370_ _2374_ _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_78_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8217__A1 as2650.stack\[4\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8217__B2 as2650.stack\[5\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8768__A2 _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6318__I _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7858__B _2744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_24_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output34_I net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_3_1_0_wb_clk_i clknet_0_wb_clk_i clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8940__A2 _3989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5754__A2 _4151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8689__B _3777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7259__A2 _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_63_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8208__A1 _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9194__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6219__B1 _4544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6228__I _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5132__I as2650.r123\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5442__A1 _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5442__B2 _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4971__I _4550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4930_ _4509_ _4510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5993__A2 _4167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7195__A1 _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4861_ _4211_ _4442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6600_ _1828_ _1829_ _1830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7580_ _1582_ _2705_ _2709_ _4268_ _2714_ _2715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_4792_ _4300_ _4372_ _4373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6531_ _1763_ _1764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9250_ _0143_ clknet_leaf_64_wb_clk_i as2650.r123\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8695__A1 _4441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6462_ _1504_ _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8201_ _2440_ _3302_ _3305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5413_ as2650.holding_reg\[6\] _0718_ _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6393_ _0985_ _1643_ _1647_ _0057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_9181_ _0074_ clknet_leaf_8_wb_clk_i as2650.ins_reg\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6170__A2 _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8132_ _2633_ _3237_ _3241_ _3242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8447__A1 _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5344_ _0418_ _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8998__A2 _4027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8063_ _2618_ _0687_ _2607_ _3176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5275_ as2650.r123\[2\]\[5\] as2650.r123_2\[2\]\[5\] _0493_ _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7522__I _2340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7014_ _2162_ _2212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8781__C _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8965_ _0846_ _3987_ _4006_ _4007_ _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5977__I _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5433__A1 _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7916_ net52 _2942_ _2943_ _3043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xclkbuf_leaf_37_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_102_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8896_ as2650.stack\[7\]\[13\] _3947_ _3956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5984__A2 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7847_ _2960_ _2975_ _2976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_51_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7778_ _0966_ _2684_ _2908_ _2681_ _2909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_51_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5736__A2 _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6729_ _1867_ _1896_ _1943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_20_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8686__A1 _4316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_9379_ _0272_ clknet_leaf_45_wb_clk_i as2650.psu\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5217__I _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8438__A1 _2495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7860__C _2661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8438__B2 _3533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8989__A2 _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7432__I _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5121__B1 _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7588__B _2722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8610__A1 _3492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6621__B1 _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8263__I _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7177__A1 _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8913__A2 _3969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5727__A2 _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6511__I _1744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8866__C _3933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8429__A1 _3379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4966__I _4545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7342__I _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5060_ _0369_ _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5663__A1 _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8601__A1 _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8750_ _0924_ _3758_ _3825_ _3835_ _3836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_92_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5962_ _4426_ _1235_ _4489_ _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__5966__A2 _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7701_ _1599_ _0830_ _2832_ _2833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_0_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4913_ _4493_ _4494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8681_ _4428_ _4137_ _3770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7168__A1 _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8365__B1 _3464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5893_ _0578_ _1096_ _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7632_ _2759_ _2765_ _2766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8901__I _3958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4844_ _4424_ _4425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_14_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7563_ _2695_ _2697_ _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_105_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4775_ as2650.addr_buff\[6\] _4355_ _4356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_9302_ _0195_ clknet_leaf_1_wb_clk_i as2650.holding_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6514_ _1745_ _1748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7494_ _2629_ _2630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9233_ _0126_ clknet_3_0_0_wb_clk_i as2650.r123_2\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6445_ _1678_ _1686_ _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7340__A1 _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5037__I as2650.r123\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9164_ _0057_ clknet_leaf_48_wb_clk_i as2650.stack\[3\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7891__A2 _3017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6376_ _1568_ _1574_ _1632_ _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8115_ _1328_ _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5327_ _0540_ _4499_ _0634_ _0004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__9093__A1 _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9095_ _4125_ _4122_ net27 _4126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_130_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8046_ _1676_ _1268_ _3159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6446__A3 _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5258_ _0542_ _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5189_ as2650.r0\[4\] _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7946__A3 _3070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8948_ _3994_ _3996_ _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5500__I _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5957__A2 _4227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7159__A1 _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8879_ _2307_ _3935_ _3945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_12_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5709__A2 _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7427__I _2564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6331__I _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8659__A1 _2927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7331__A1 _2469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7882__A2 _2522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5893__A1 _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9084__A1 _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7162__I _2315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7634__A2 _2686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8831__A1 _2285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5645__A1 _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5611__S _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9232__CLK clknet_leaf_63_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6070__A1 _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9382__CLK clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9038__B _3868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7570__A1 _2565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4560_ _4140_ _4141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7322__A1 _4161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8665__A4 _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6230_ _1486_ _1487_ _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_83_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5884__A1 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4696__I _4192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6161_ as2650.stack\[4\]\[11\] _1420_ _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__9075__A1 _4100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7072__I _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5112_ _0421_ _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6092_ _1282_ _1362_ _1363_ _1364_ _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__7625__A2 _2749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5636__A1 _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5043_ _0352_ _0287_ _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5100__A3 _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8117__B _3207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7928__A3 _3052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6416__I _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8802_ _0944_ _3856_ _3245_ _3885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6994_ _2194_ _2195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5939__A2 _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6061__A1 _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8733_ _3763_ _3808_ _3809_ _3819_ _3820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_129_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5945_ _0830_ _1059_ _1136_ _1219_ _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_55_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8664_ _3752_ _3753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8889__A1 _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6349__C1 _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5876_ _0446_ _0474_ _1082_ _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_90_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7615_ _2748_ _2749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4827_ _4154_ _4407_ _4408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8595_ _0995_ _0988_ _3648_ _3687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7546_ _2183_ _2580_ _2680_ _2681_ _2682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4758_ _4330_ _4335_ _4336_ _4337_ _4338_ _4339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_120_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4914__A3 _4486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7477_ _2606_ _2608_ _2611_ _2613_ _2570_ _2614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__6116__A2 _4527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7313__A1 _2450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4689_ _4247_ _4262_ _4269_ _4270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_49_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9216_ _0109_ clknet_leaf_41_wb_clk_i as2650.stack\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6428_ _1011_ _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5875__A1 _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4678__A2 _4257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9147_ _0040_ clknet_leaf_15_wb_clk_i net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9066__A1 _4100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6359_ net3 _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7616__A2 _2746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9078_ _3132_ _4105_ _4111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9255__CLK clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_52_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_52_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_8029_ _1706_ _1572_ _3145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4850__A2 _4313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6052__A1 _4174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7866__B _2483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6996__I _2196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7304__A1 _1497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9057__A1 _3851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6010__B _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8804__A1 _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7620__I _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7776__B _2624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7791__A1 _2919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6594__A2 _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5730_ _0959_ _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5661_ _0850_ _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7543__A1 _2658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6346__A2 _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7400_ _2154_ _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9128__CLK clknet_leaf_58_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4612_ _4158_ _4177_ _4193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8380_ _3458_ _3457_ _3479_ _3291_ _3480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_5592_ _0895_ _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_50_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7331_ _2469_ _4352_ _2470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7262_ _4323_ _2401_ _2402_ _1410_ _0171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__7846__A2 _2974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5857__A1 _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9001_ _4479_ _0624_ _4040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__9048__A1 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6213_ _4255_ _4232_ _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_7193_ _0852_ _1283_ _4253_ _2343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_63_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6144_ _1397_ _1408_ _1409_ _1410_ _0045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6075_ _4164_ _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5085__A2 _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6282__A1 _4328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5026_ _4542_ _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4832__A2 _4353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8023__A2 _3103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5050__I _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6977_ _2179_ _2180_ _0108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8716_ _3703_ _3803_ _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5928_ _1056_ _1201_ _1203_ _1053_ _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__5918__C _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8326__A3 _3355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8647_ _3724_ _3148_ _3736_ _3194_ _3737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7534__A1 _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5859_ _0422_ _1094_ _1138_ _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_107_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8578_ _3392_ _3665_ _3671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4899__A2 _4479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7529_ _2663_ _2664_ _2665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5848__A1 _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9039__A1 _3088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8262__A2 _3361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7440__I _2577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_40_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6273__A1 _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4823__A2 _4377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6056__I _4235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8014__A2 _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6025__A1 _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7773__A1 _2884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5379__A3 _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8271__I _3373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7525__A1 _2336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5839__A1 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8253__A2 _3301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6264__A1 _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5067__A2 _4507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4814__A2 _4393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6900_ _2005_ _2109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7880_ _1546_ _3006_ _3007_ _2852_ _3008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_75_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6016__A1 _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6831_ _2033_ _2042_ _2043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_90_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6762_ _1952_ _1975_ _1976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_108_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8501_ as2650.pc\[8\] _2203_ _3570_ _3597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_5713_ _1003_ _0980_ _0972_ as2650.r123_2\[0\]\[4\] _1004_ _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_91_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7516__A1 _2648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6693_ as2650.stack\[1\]\[13\] _1907_ _1916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7516__B2 _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8432_ _0946_ _3529_ _3530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_104_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5644_ _0915_ _0942_ _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8363_ _2188_ _1605_ _3463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5575_ _0878_ _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7314_ _2406_ _2448_ _2452_ _2453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7819__A2 _2876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8294_ _0920_ _3355_ _3396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_116_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7245_ _1466_ _2387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7176_ _2302_ _2313_ _2316_ as2650.stack\[0\]\[5\] _2310_ _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_59_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6127_ _1373_ _1395_ _1396_ _1392_ _0042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8244__A2 _2438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5058__A2 _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6058_ _1328_ _1330_ _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_14_wb_clk_i_I clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4805__A2 _4385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5009_ _0300_ _0319_ _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6007__A1 _4430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7755__A1 _2884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8305__B _3406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8952__B1 _3993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5230__A2 _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7435__I _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4741__A1 _4321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8483__A2 _3569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_53_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5297__A2 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4794__I _4374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8266__I _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8235__A2 _3335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6246__A1 _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7994__A1 _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8538__A3 _3632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7746__A1 _1604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6549__A2 _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6514__I _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5221__A2 _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8869__C _3933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4980__A1 _4348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4980__B2 _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8171__A1 _2439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7345__I _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6721__A2 _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4732__A1 _4159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5360_ _0610_ _0590_ _0663_ _4350_ _0666_ _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_114_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8474__A2 _3570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5291_ _4508_ _0480_ _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7030_ _2178_ _2219_ _2220_ as2650.stack\[4\]\[2\] _2221_ _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_101_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6237__A1 _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7434__B1 _2567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9316__CLK clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8981_ _3057_ _0897_ _2408_ _1272_ _4021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_55_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6788__A2 _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7932_ _3057_ _3058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8904__I _3961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5460__A2 _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7863_ _0989_ _0757_ _2991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7737__A1 _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6814_ _1996_ _2024_ _2025_ _2026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5468__C _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7794_ _2818_ _2915_ _2922_ _2923_ _2924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5212__A2 _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6745_ _1843_ _1884_ _1959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6960__A2 _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6676_ _1903_ _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8162__A1 _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8415_ _3059_ _3503_ _3510_ _3513_ _3514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5627_ _0927_ _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8346_ as2650.stack\[3\]\[3\] _1919_ _1638_ as2650.stack\[2\]\[3\] _3447_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_5558_ as2650.pc\[0\] _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8465__A2 _3561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8277_ _3291_ _3379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5489_ as2650.holding_reg\[7\] _4376_ _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_120_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7228_ _2373_ _2359_ _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4828__B _4408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7159_ _2146_ _2313_ _2316_ as2650.stack\[0\]\[0\] _2310_ _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__8217__A2 _3319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7976__A1 _1692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output27_I net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7728__A1 _2204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6400__A1 as2650.stack\[3\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8153__A1 _2484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7900__A1 net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8456__A2 _3366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6467__A1 _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__9339__CLK clknet_leaf_51_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8208__A2 _2854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6219__A1 _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6219__B2 _4199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7967__A1 _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5442__A2 _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7719__A1 _2491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4860_ _4406_ _4441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7195__A2 _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4791_ as2650.r123\[1\]\[7\] as2650.r123\[0\]\[7\] as2650.r123_2\[1\]\[7\] as2650.r123_2\[0\]\[7\]
+ _4197_ _4148_ _4372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6530_ _1762_ _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4953__A1 _4249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8144__A1 _2150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6461_ _1700_ _0072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_88_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8200_ _2145_ _3302_ _3303_ _3304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4705__A1 _4138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5412_ _0717_ _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_127_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9180_ _0073_ clknet_leaf_6_wb_clk_i as2650.ins_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6392_ as2650.stack\[3\]\[9\] _1646_ _1647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6170__A3 _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8131_ _3239_ _3240_ _4201_ _3241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5343_ _0555_ _0648_ _0649_ _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_114_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8062_ _4241_ _3175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5274_ _4521_ _0581_ _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7013_ _2210_ _2211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6419__I _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7958__A1 _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8634__I as2650.pc\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8964_ _2131_ _2132_ _2135_ _3962_ _4007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__6630__A1 _1795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5433__A2 _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5479__B _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7915_ _1003_ _2522_ _3041_ _2940_ _3042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_37_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8895_ _1670_ _3949_ _3955_ _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8907__B1 _3964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5984__A3 _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7846_ _2961_ _2974_ _2975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_77_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_77_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_75_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7777_ _2889_ _2898_ _2906_ _2907_ _2908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_71_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4989_ _4279_ _0299_ _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6728_ _1941_ _1942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4944__A1 _4518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8135__A1 _1486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4830__C _4345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6659_ _0364_ _1887_ _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8686__A2 _3772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9378_ _0271_ clknet_leaf_8_wb_clk_i as2650.ins_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_139_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8329_ _1293_ _3353_ _3430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5121__A1 as2650.stack\[0\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8610__A2 _3686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6621__A1 _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6621__B2 _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8374__A1 as2650.addr_buff\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6999__I _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6924__A2 _2114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8126__A1 _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6688__A1 _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9161__CLK clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8429__A2 _3495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5360__A1 _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5360__B2 _4350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7623__I net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6239__I _4255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5663__A2 _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8601__A2 _2776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6612__A1 as2650.r0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5961_ _4433_ _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_3_2_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7700_ _2806_ _2809_ _2831_ _2832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4912_ _4415_ _4492_ _4493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8680_ _1235_ _3769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5892_ _0500_ _1063_ _1169_ _1058_ _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__8365__A1 _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8365__B2 _2524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7631_ _2499_ _2763_ _2764_ _2765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5179__A1 _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4843_ _4312_ _4423_ _4424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6915__A2 _2114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6702__I _1922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7562_ _2636_ _2696_ _2697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__8117__A1 _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4774_ as2650.addr_buff\[5\] _4355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_144_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9301_ _0194_ clknet_leaf_1_wb_clk_i as2650.holding_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6513_ _4284_ _1746_ _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7493_ _1283_ _2629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8668__A2 _3750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5318__I _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9232_ _0125_ clknet_leaf_63_wb_clk_i as2650.r123_2\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6444_ _1680_ _1685_ _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7340__A2 _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9163_ _0056_ clknet_leaf_48_wb_clk_i as2650.stack\[3\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6375_ _1576_ _1548_ _1631_ _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_66_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8114_ _3210_ _3218_ _3224_ _3225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5326_ _4500_ _0616_ _0633_ _0538_ _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_138_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9094_ _1588_ _4113_ _4125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9093__A2 _4113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8045_ _3157_ _3158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5257_ _0562_ _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6446__A4 _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5053__I _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5188_ _4298_ _0496_ _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7800__B1 _2688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8947_ _3995_ _2017_ _3996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8356__A1 _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8878_ _2305_ _3931_ _3932_ as2650.stack\[7\]\[7\] _3923_ _3944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7829_ _2613_ _2947_ _2957_ _2888_ _2958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_58_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6906__A2 _2114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9184__CLK clknet_leaf_69_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5590__A1 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8659__A2 _3747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7871__C _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7331__A2 _4352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7443__I _2517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5893__A2 _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9084__A2 _3136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8831__A2 _3908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8274__I _3376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8595__A1 _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6070__A2 _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8347__A1 as2650.stack\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8898__A2 _3947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4908__A1 _4143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7570__A2 _2704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5138__I _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7322__A2 _2458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9054__B _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5333__A1 _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7353__I _2491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6160_ _0993_ _1417_ _1422_ _0049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_112_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5111_ _0396_ _0419_ _0420_ _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7086__A1 _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6091_ _1315_ _0882_ _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5042_ _4349_ _4244_ _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_57_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8184__I _3287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8801_ _2458_ _2753_ _3877_ _3883_ _3884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7928__A4 _3053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6993_ as2650.pc\[5\] _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_19_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6061__A2 _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8912__I _3958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5944_ _1058_ _1218_ _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8732_ _1699_ _3766_ _2629_ _3818_ _3819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_94_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8663_ _4242_ _2469_ _1491_ _3751_ _3752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_55_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6349__B1 _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8889__A2 _3948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5875_ _0485_ _1134_ _1152_ _1153_ _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6349__C2 _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7010__A1 _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7614_ net33 _2747_ _2748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_107_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4826_ _4157_ _4268_ _4407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8594_ _3685_ _3686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7545_ _2403_ _2681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4757_ _4226_ _4338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4914__A4 _4494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7476_ _2612_ _2613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4688_ _4233_ _4206_ _4268_ _4269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_88_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8510__A1 _3533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7313__A2 _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8359__I _3394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6427_ _1670_ _1661_ _1671_ _0067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_9215_ _0108_ clknet_leaf_41_wb_clk_i as2650.stack\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7263__I _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9146_ _0039_ clknet_leaf_15_wb_clk_i net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5875__A2 _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4678__A3 _4245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6358_ _1593_ _1610_ _1613_ _1614_ _1615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_115_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5309_ _0580_ _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9077_ _4107_ _4110_ _3619_ _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8813__A2 _3894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6289_ _1540_ _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8028_ _3143_ _3144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8329__A1 _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8501__A1 as2650.pc\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7304__A2 _4250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9057__A2 _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6010__C _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7607__A3 _2707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8804__A2 _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8568__A1 _3379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8568__B2 _3661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5660_ _0956_ _0015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7543__A2 _2660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4611_ _4183_ _4192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_129_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5591_ _0884_ _4208_ _0894_ _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_50_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7330_ _2468_ _2469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7261_ net22 _2401_ _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9000_ _3492_ _3122_ _4026_ _4039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5857__A2 _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6212_ _4543_ _1361_ _1470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_144_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7192_ _2150_ _1532_ _0871_ _2342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__9048__A2 _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6143_ _1391_ _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6074_ _1346_ _4237_ _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5025_ _4485_ _0335_ _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8559__A1 _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7967__B _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6034__A2 _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6976_ _0918_ _2176_ _2180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7782__A2 _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8715_ _1382_ _3758_ _3802_ _3803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5927_ _0783_ _1117_ _1202_ _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__5793__A1 _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7258__I _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8031__I0 _3146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8646_ _2634_ _3727_ _3736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_16_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5858_ _1132_ _1135_ _1137_ _1094_ _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_107_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8731__A1 _3767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8798__B _3880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4809_ net6 _4390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8577_ _3668_ _3669_ _3670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5789_ _1070_ _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7528_ _1584_ _0479_ _0484_ _2664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_108_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8310__C _3411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7298__A1 _1497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7459_ _1553_ _2592_ _2595_ _2596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__9222__CLK clknet_leaf_40_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5848__A2 _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9039__A2 _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9129_ _0022_ clknet_leaf_58_wb_clk_i as2650.stack\[6\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8798__A1 _1627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9372__CLK clknet_leaf_76_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6273__A2 _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6337__I _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7773__A2 _2618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5379__A4 _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8970__A1 _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7525__A2 _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8722__A1 _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7289__A1 _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8486__B1 _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5839__A2 _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8789__A1 _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6264__A2 _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5472__B1 _4469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4814__A3 _4394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6016__A2 _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6830_ _2001_ _2041_ _2042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_1_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8961__A1 _3966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6761_ _1958_ _1974_ _1975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_62_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7078__I _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8500_ _3595_ _3596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5712_ _0540_ _4416_ _0982_ _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6692_ _1670_ _1909_ _1915_ _0088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_56_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7516__A2 _2650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8713__A1 _3088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8431_ _2195_ _3494_ _3529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5643_ _0940_ _0904_ _0941_ _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__9245__CLK clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8411__B _3504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8362_ _3460_ _3461_ _1685_ _3462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5574_ _4207_ _4175_ _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7313_ _2450_ _1503_ _2451_ _2452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_116_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8293_ _3394_ _3395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7819__A3 _2878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7244_ _2385_ _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7175_ _0932_ _2311_ _2328_ _0158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_67_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6126_ net44 _1380_ _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_24_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7452__A1 _2584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6057_ _1329_ _1306_ _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5061__I _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5008_ _4338_ _0303_ _0317_ _0318_ _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_73_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6007__A2 _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7755__A2 _2885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8952__A1 _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5766__A1 _4195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6959_ _0900_ _2165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8004__I0 _3124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5518__A1 _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5945__B _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8629_ _0709_ _3481_ _3426_ _3706_ _3719_ _3720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__5369__I1 as2650.r123\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6191__A1 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5236__I _4325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4741__A2 _4311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7691__A1 _2774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7451__I _4246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6067__I _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6246__A2 _4550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__9118__CLK clknet_leaf_39_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7994__A2 _2420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7746__A2 _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9268__CLK clknet_leaf_52_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_7_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5855__B _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8171__A2 _3186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6182__A1 _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4732__A2 _4179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5390__C1 _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5290_ _4396_ _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4985__I _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7682__A1 _2729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7361__I _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7434__A1 _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6237__A2 _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7434__B2 _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8980_ _2342_ _2400_ _4016_ _4019_ _4020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_110_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7985__A2 _3107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7931_ _2157_ _3057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5996__A1 _4201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7862_ as2650.pc\[11\] _1586_ _2990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_110_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7737__A2 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8934__A1 _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6813_ _1999_ _2012_ _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5748__A1 as2650.stack\[5\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7793_ _2570_ _2923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6744_ _1956_ _1957_ _1958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_52_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6675_ _1902_ _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8162__A2 _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5626_ _0926_ _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8414_ _3395_ _3511_ _3512_ _3513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_104_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8345_ _3445_ _3446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5920__A1 _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5557_ _0860_ _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8276_ _3375_ _3378_ _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5488_ _0787_ _0792_ _4498_ _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_65_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7673__A1 _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4895__I _4475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7227_ _1558_ _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7158_ _2315_ _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6109_ _1373_ _1379_ _1381_ _1302_ _0039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_112_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5005__B _4324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8622__B1 _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7089_ _0947_ _2265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7728__A2 _2496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5739__A1 _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8830__I _3900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8153__A2 _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5394__C _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6164__A1 _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5911__A1 _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9102__A1 _3132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7664__A1 _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8277__I _3291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6219__A2 _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5630__S _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8226__B _3329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7719__A2 _2646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8916__A1 _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_33_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4790_ _4369_ _4370_ _4371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4953__A2 _4258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7356__I _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8144__A2 _3250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6260__I _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6460_ _1696_ _1688_ _1698_ _1699_ _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6155__A1 _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_12_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5411_ _0716_ _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4705__A2 _4135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6391_ _1641_ _1646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8130_ _2624_ _3061_ _1339_ _2390_ _3240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_127_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5342_ _0640_ _0647_ _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_114_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8187__I _3290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8061_ _1677_ _3153_ _2407_ _3173_ _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_99_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5273_ as2650.r123\[1\]\[5\] as2650.r123\[0\]\[5\] as2650.r123_2\[1\]\[5\] as2650.r123_2\[0\]\[5\]
+ _4196_ _0493_ _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_88_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7012_ _2209_ _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5130__A2 _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7958__A2 _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8963_ as2650.r123\[2\]\[7\] _3989_ _4006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6435__I _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7914_ _3018_ _3019_ _3034_ _3040_ _3041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__6630__A2 _1859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8894_ as2650.stack\[7\]\[12\] _3951_ _3955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8907__A1 _3962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8907__B2 as2650.r123\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7845_ _2934_ _2912_ _2974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_54_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8383__A2 _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7776_ _0966_ _2528_ _2624_ _2907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4988_ _0297_ _4332_ _0298_ _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6727_ _1939_ _1035_ _1940_ _4438_ _1941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__7266__I _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4944__A2 _4523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8135__A2 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6146__A1 _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6658_ _1781_ _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5609_ _0911_ _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_46_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_46_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6697__A2 _4458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9377_ _0270_ clknet_leaf_9_wb_clk_i as2650.ins_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6589_ _1814_ _1819_ _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_69_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8328_ _0920_ _3355_ _2182_ _3429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_11_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7646__A1 _2757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8097__I _3207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8259_ _1655_ _3362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5121__A2 _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8825__I _3905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4632__A1 _4195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8374__A2 _2754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5188__A2 _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8126__A2 _2506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6137__A1 _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7885__A1 as2650.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6688__A2 _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4699__A1 _4138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5852__C _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6255__I _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5960_ _4443_ _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4623__A1 _4201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4911_ _4436_ _4491_ _4492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5891_ _1076_ _1168_ _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8365__A2 _3457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7630_ _2757_ _1614_ _2764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5179__A2 _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4842_ _4224_ _4278_ _4423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7561_ _2601_ _2619_ _2637_ _2639_ _2696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4773_ _4269_ _4354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8117__A2 _3227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9300_ _0193_ clknet_leaf_1_wb_clk_i as2650.holding_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6512_ _1745_ _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7492_ _2579_ _2627_ _2628_ _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8668__A3 _3755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9231_ _0124_ clknet_leaf_61_wb_clk_i as2650.r123_2\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6443_ _1684_ _1685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7340__A3 _4240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9162_ _0055_ clknet_leaf_45_wb_clk_i as2650.psl\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6374_ _1577_ _1630_ _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7628__A1 _2727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8113_ _3220_ _3222_ _3223_ _3224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5325_ _0617_ _0621_ _4446_ _0632_ _0438_ _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_66_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9093_ _0944_ _4113_ _4123_ _4124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8044_ _2503_ _3157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5256_ _0554_ _0563_ _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5187_ as2650.r123\[2\]\[4\] as2650.r123_2\[2\]\[4\] _4516_ _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_56_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8053__A1 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7800__A1 _2919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7800__B2 _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8946_ _3961_ _3995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4614__A1 _4191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8877_ _2199_ _3925_ _3943_ _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8356__A2 _3455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7828_ _2951_ _2956_ _2661_ _2957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__9329__CLK clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7759_ as2650.pc\[8\] _0755_ _2890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_36_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5509__I _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7724__I _2855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5342__A2 _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9084__A3 _4100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8292__A1 _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4853__A1 _4426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4605__A1 _4179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6358__A1 _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6358__B2 _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4908__A2 _4488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5030__A1 _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6024__B _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7322__A3 _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5333__A2 _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5110_ _0395_ _0408_ _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6090_ _4550_ _0879_ _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8283__B2 as2650.stack\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5041_ _0348_ _0350_ _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_0_wb_clk_i wb_clk_i clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_8800_ _1588_ _3766_ _3881_ _3882_ _2630_ _3883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_80_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6992_ _0937_ _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8731_ _3767_ _1393_ _3817_ _3765_ _3818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_80_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5943_ _0789_ _1110_ _1217_ _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_59_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8662_ _1328_ _1338_ _1496_ _2448_ _3751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__6349__A1 _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7546__B1 _2680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5874_ _0491_ _1097_ _1134_ _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6349__B2 _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8133__C _3229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7613_ net32 _2690_ _2747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_22_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7010__A2 _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4825_ _4405_ _4406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8593_ _3035_ _3684_ _3685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5329__I _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7544_ _0928_ _2630_ _2633_ _2657_ _2679_ _2680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__7972__C _2525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4756_ _4290_ _4293_ _4337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_119_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7849__A1 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7475_ _1306_ _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4687_ _4263_ _4267_ _4268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_134_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7313__A3 _2451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9214_ _0107_ clknet_leaf_41_wb_clk_i as2650.stack\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6426_ as2650.stack\[2\]\[12\] _1664_ _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6521__A1 _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5324__A2 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4678__A4 _4258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9145_ _0038_ clknet_leaf_6_wb_clk_i as2650.psu\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5064__I _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6357_ _0837_ _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5308_ _4276_ _0570_ _0609_ _0615_ _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_62_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6288_ _1545_ _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9076_ _3138_ _4108_ _4109_ _4110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5088__A1 as2650.holding_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5999__I _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8027_ _1524_ _3143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5239_ _0543_ _0546_ _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_40_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8577__A2 _3669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9151__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8929_ as2650.r123\[1\]\[6\] _3967_ _3980_ _3981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_38_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5260__A1 _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8329__A2 _3353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_61_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_61_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_130_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8501__A2 _2203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5315__A2 _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8265__A1 _3360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9321__D _0214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5702__I as2650.pc\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4826__A1 _4157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8017__A1 _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5251__A1 _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8740__A2 _3451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4610_ _4190_ _4191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7792__C _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5590_ _0893_ _4164_ _4172_ _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7364__I _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6503__A1 _1735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7260_ _2399_ _1278_ _1242_ _2400_ _2401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_144_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6211_ _0340_ _1468_ _1429_ _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7191_ _1317_ _2340_ _1496_ _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6142_ net20 _1402_ _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_139_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6073_ _4167_ _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_97_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5612__I _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9174__CLK clknet_leaf_60_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5024_ _0325_ _0330_ _0334_ _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__8008__A1 _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8559__A2 _3406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7231__A2 _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8144__B _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6975_ _2178_ _2171_ _2172_ as2650.stack\[2\]\[2\] _2173_ _2179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__6443__I _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8714_ _3763_ _3788_ _3801_ _3802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5926_ _0781_ _1119_ _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6990__A1 _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8645_ _3728_ _3734_ _3293_ _3735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5857_ _0358_ _1136_ _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8731__A2 _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8798__C _3851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4808_ _4229_ _4389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8576_ _2998_ _2538_ _3021_ _3609_ _3669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5788_ _4395_ _1037_ _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4898__I _4478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7527_ _1585_ _0485_ _2663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_135_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4739_ as2650.psl\[3\] _4320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7298__A2 _4543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7207__C _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7458_ _2593_ _2561_ _2594_ _2595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6409_ _0851_ _1657_ _0960_ _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_7389_ _2526_ _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8247__A1 _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5950__C _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9128_ _0021_ clknet_leaf_58_wb_clk_i as2650.stack\[6\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8798__A2 _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9059_ _4316_ _4078_ _4094_ _3742_ _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_89_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5233__A1 _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8970__A2 _2634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6981__A1 _2183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8722__A2 _2632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5536__A2 _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9316__D _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4601__I as2650.ins_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8486__A1 as2650.stack\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7289__A2 _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9197__CLK clknet_leaf_47_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8238__A1 _4530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8789__A2 _3856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8410__A1 _2509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5224__A1 _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8961__A2 _2129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6760_ _1960_ _1973_ _1974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_51_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6972__A1 _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5711_ _1002_ _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6691_ as2650.stack\[1\]\[12\] _1911_ _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8430_ _0940_ _3289_ _3528_ _3112_ _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_104_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5642_ as2650.stack\[5\]\[5\] _0913_ _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8411__C _3509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8361_ _2189_ _3428_ _3461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_141_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5573_ _0876_ _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5607__I _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7312_ _4220_ _2406_ _0970_ _2451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8477__A1 _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8292_ _1271_ _2157_ _3155_ _3394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_85_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7243_ _2384_ _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8229__A1 _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7174_ _2300_ _2313_ _2316_ as2650.stack\[0\]\[4\] _2310_ _2328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_113_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6438__I _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6125_ _0924_ _1376_ _1394_ _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_100_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6056_ _4235_ _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5463__A1 _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5007_ _4330_ _0304_ _4338_ _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_73_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8401__A1 _4265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8952__A2 _3992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5766__A2 _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6963__A1 _2147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6958_ _2163_ _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6963__B2 as2650.stack\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5909_ _0698_ _1096_ _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8004__I1 _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6889_ _2073_ _2098_ _2099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_70_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8628_ _3715_ _3717_ _3718_ _3719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5945__C _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6715__A1 _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8180__A3 _3283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8559_ _2395_ _3406_ _3653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6191__A2 _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8468__A1 _2825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8828__I _3903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7140__A1 _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6348__I _1604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7888__B _2825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8640__A1 as2650.pc\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5454__A1 _4533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5057__I1 as2650.r123\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6083__I _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5757__A2 _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8004__S _3120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6706__A1 _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5390__C2 _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5871__B _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7131__A1 _2294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7682__A2 _2727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5693__A1 _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6258__I _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7434__A2 _2537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8631__A1 _3379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7930_ _3044_ _2462_ _3054_ _3055_ _3056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_110_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5996__A2 _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7861_ _2613_ _2984_ _2988_ _2888_ _2989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7089__I _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8934__A2 _3959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6812_ _1999_ _2012_ _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7792_ _2836_ _2918_ _2921_ _2720_ _2486_ _2922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__6945__A1 _2150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5748__A2 _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6743_ _0499_ _1887_ _1957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9362__CLK clknet_leaf_69_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6674_ _4467_ _4457_ _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8413_ _0940_ _3460_ _3512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5625_ as2650.pc\[3\] _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6173__A2 _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4803__S0 _4139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8344_ _3415_ _3424_ _3433_ _2524_ _2856_ _3445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5556_ _0859_ _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_3_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8275_ _2170_ _3377_ _1566_ _3378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5487_ _0791_ _0620_ _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_133_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7226_ as2650.addr_buff\[4\] _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__7673__A2 _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8870__A1 _2298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7157_ _2165_ _2314_ _2315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6108_ net41 _1380_ _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8622__A1 _4265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8622__B2 _3712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7088_ _2193_ _2245_ _2264_ _0135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_98_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6484__I0 as2650.r123\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6039_ _1309_ _1310_ _1311_ _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_73_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5800__I _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7189__A1 _2335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8925__A2 _3967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5739__A2 _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8689__A1 _3768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5247__I _4315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5911__A2 _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9102__A2 _4121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8310__B1 _3409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5124__B1 _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7664__A2 _2686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9235__CLK clknet_leaf_62_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8293__I _3394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5710__I as2650.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8916__A2 _3969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6927__A1 _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8129__B1 _3178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7637__I _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7352__A1 _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5410_ _0673_ _0675_ _0677_ _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_51_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6390_ _0976_ _1643_ _1645_ _0056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_103_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5341_ _0641_ _0647_ _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8060_ _3154_ _3161_ _3165_ _3172_ _3173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_5272_ _0579_ _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_99_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5106__B _4314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7011_ _1018_ _2208_ _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7958__A3 _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8962_ _4004_ _4005_ _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5969__A2 _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6091__A1 _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7913_ _1450_ _3039_ _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_fanout51_I net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7040__C _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8893_ _1668_ _3948_ _3954_ _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_3_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7844_ _0990_ _2513_ _2972_ _2928_ _2551_ _2973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_52_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7040__B1 _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7775_ _2901_ _2905_ _2550_ _2906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8152__B _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7591__A1 _2579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4987_ _4257_ _4386_ _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6726_ _1612_ _1051_ _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_71_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8135__A3 _3209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6657_ _1874_ _1879_ _1885_ _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__6146__A2 _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5608_ _0910_ _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__9108__CLK clknet_leaf_68_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7894__A2 as2650.addr_buff\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9376_ _0269_ clknet_leaf_74_wb_clk_i as2650.r123\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6588_ _1815_ _1817_ _1818_ _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_139_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8327_ _3427_ _3428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5539_ _0790_ _4547_ _0842_ _0843_ _0486_ _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_117_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8258_ _1903_ _3361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8843__A1 _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5657__A1 as2650.stack\[5\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9258__CLK clknet_leaf_56_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7209_ _2357_ _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_15_wb_clk_i clknet_3_2_0_wb_clk_i clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_132_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8189_ _3095_ _3293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5530__I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9002__I _3122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4632__A2 _4212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9020__A1 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6909__B2 _1980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7582__A1 _2636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6385__A2 _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6361__I _1617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7885__A2 _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8598__B1 _3689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4910_ _4490_ _4491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__9011__A1 _4026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5890_ _0371_ _1127_ _1167_ _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4841_ _4421_ _4422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_60_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6376__A2 _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7560_ _2187_ _2694_ _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4772_ _4352_ _4353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_140_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6511_ _1744_ _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7491_ _2609_ _2466_ _1635_ _2628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8668__A4 _3756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9230_ _0123_ clknet_leaf_61_wb_clk_i as2650.r123_2\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6442_ _1683_ _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_23_wb_clk_i_I clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5887__A1 _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9161_ _0054_ clknet_3_4_0_wb_clk_i as2650.psl\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__9078__A1 _3132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6373_ _1621_ _1625_ _1626_ _1627_ _1629_ _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__6220__B _4419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_3_0_0_wb_clk_i clknet_0_wb_clk_i clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__5615__I _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8112_ _4253_ _3153_ _2508_ _3059_ _3191_ _3223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_114_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5324_ _0628_ _0631_ _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9092_ _1706_ _4028_ _4123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8043_ _1250_ _3155_ _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5255_ _0555_ _0558_ _0561_ _0418_ _0562_ _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_87_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5186_ _4521_ _0494_ _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8053__A2 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7800__A2 _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8945_ _0323_ _3992_ _3993_ as2650.r123\[2\]\[1\] _3994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4614__A2 _4194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8876_ _0948_ _3927_ _3929_ as2650.stack\[7\]\[6\] _3933_ _3943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_97_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7827_ _2954_ _2955_ _2366_ _2956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7277__I _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_62_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7758_ _2836_ _2883_ _2887_ _2888_ _2889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_51_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6709_ _1663_ _1924_ _1928_ _0092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_71_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7316__A1 _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7689_ _2201_ _2684_ _2821_ _2681_ _2822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__8610__B _3331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5590__A3 _4172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9069__A1 _2793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9359_ _0252_ clknet_leaf_59_wb_clk_i as2650.stack\[7\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5525__I _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8816__A1 _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7740__I _2867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8292__A2 _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6055__A1 _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8595__A3 _3648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9319__D _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4908__A3 _4432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6024__C _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5030__A2 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7307__A1 _4422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7858__A2 _2950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5869__A1 _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8807__A1 _3838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8283__A2 _3319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5040_ _0349_ _4509_ _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6266__I _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6991_ _2186_ _2143_ _2192_ _0110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_65_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7794__A1 _2818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8730_ _3790_ _3816_ _3817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5942_ _0680_ _1127_ _1214_ _1216_ _1062_ _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_111_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8661_ _1463_ _3748_ _3749_ _3265_ _3750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__7546__A1 _2183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5873_ _0535_ _1099_ _1151_ _1061_ _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_59_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6349__A2 _4334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7546__B2 _2681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7612_ _2738_ _2745_ _2746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4824_ _4285_ _4405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8592_ as2650.pc\[11\] _3663_ _3684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5021__A2 _4460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7543_ _2658_ _2660_ _2678_ _2483_ _2679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_119_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4755_ _4324_ _4336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7474_ _2609_ _2610_ _2611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7849__A2 _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4686_ as2650.addr_buff\[7\] _4266_ _4267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9213_ _0106_ clknet_leaf_56_wb_clk_i as2650.stack\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6425_ _1005_ _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6521__A2 _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9144_ _0037_ clknet_leaf_66_wb_clk_i as2650.r123_2\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_115_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6356_ _1611_ _1612_ _1264_ _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_118_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5307_ _4346_ _0614_ _4412_ _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9075_ _4100_ _3135_ _4109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6287_ _1544_ _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5088__A2 _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8026_ _3142_ _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5238_ _0443_ _0459_ _0545_ _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5169_ _4304_ _4386_ _4524_ _0463_ _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__6037__A1 _4254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6109__C _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8928_ _3976_ _1859_ _3980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8859_ _3926_ _3931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4771__A1 _4304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8501__A3 _3570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_30_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_30_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_84_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5720__B1 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7470__I _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6276__A1 _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4826__A2 _4268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8017__A2 _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7776__A1 _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5858__C _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7528__A1 _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5539__B1 _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6200__A1 _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5874__B _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7645__I net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4762__A1 _4279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6210_ _0393_ _4431_ _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_7190_ _1338_ _2340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__9081__B _3133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6141_ _0944_ _1398_ _1407_ _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8256__A2 _3343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9319__CLK clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6072_ _1307_ _1344_ _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4817__A2 _4333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5023_ _0331_ _0332_ _0333_ _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_61_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8008__A2 _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_22_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7767__A1 _2895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6974_ _0920_ _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8144__C _3178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5925_ _0740_ _1083_ _1199_ _1200_ _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_0_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8713_ _3088_ _3800_ _3801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7519__A1 _2335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8644_ _3393_ _3727_ _3733_ _3598_ _3734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_94_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7983__C _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5856_ _1041_ _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4807_ _4387_ _4388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8575_ _2950_ _3610_ _2369_ _3668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5787_ _1065_ _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7526_ _1308_ _2662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4738_ _4315_ _4318_ _4319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7457_ _4528_ _4511_ _4512_ _2594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_120_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4669_ _4249_ _4250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6408_ _1656_ _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7388_ _1695_ _2395_ _2526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9127_ _0020_ clknet_leaf_58_wb_clk_i as2650.stack\[6\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8247__A2 _1618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6339_ _4316_ _4391_ _0683_ _1595_ _1596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_88_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8319__C _3420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7455__B1 _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9058_ _4089_ _4090_ _4093_ _1576_ _4078_ _4094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_118_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8009_ _3127_ _3128_ _3129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7758__A1 _2836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8335__B _3076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8955__B1 _3989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6430__A1 _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6981__A2 _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8183__A1 _3055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4744__A1 _4192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8486__A2 _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8238__A2 _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9332__D _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6249__A1 _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8229__C _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5472__A2 _4465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7749__A1 _2876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8245__B _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8410__A2 _3508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6421__A1 _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6972__A2 _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5710_ as2650.pc\[12\] _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6690_ _1668_ _1908_ _1914_ _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8174__A1 _2631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5641_ _0939_ _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7375__I _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7921__A1 _3045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8360_ _2189_ _3428_ _3460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5572_ _4180_ _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7311_ _4442_ _2449_ _2450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_89_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8477__A2 _2849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8291_ _3392_ _3393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6488__A1 _4405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7242_ _1489_ _2384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8200__S _3303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9141__CLK clknet_leaf_67_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8229__A2 _3289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7173_ _2326_ _2327_ _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5623__I _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6124_ _1377_ _1393_ _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9291__CLK clknet_leaf_31_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6055_ _1316_ _1327_ _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7978__C _2578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6660__A1 _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5006_ _0309_ _0312_ _0313_ _0316_ _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__6660__B2 _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8401__A2 _3157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6957_ _2148_ _1657_ _2162_ _2163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_74_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5908_ _0670_ _1063_ _1184_ _1058_ _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6888_ _2021_ _2047_ _2074_ _2050_ _2098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_35_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8165__A1 _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8602__C _3676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8627_ _3257_ _3706_ _3712_ _2549_ _2856_ _3718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5839_ _0335_ _1119_ _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7912__A1 _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7912__B2 _3001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5369__I3 as2650.r123_2\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4702__I _4282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8558_ _0989_ _3644_ _3652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_108_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6122__C _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6191__A3 _1428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7509_ _2352_ _2645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8468__A2 _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8489_ _3585_ _3586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_135_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6403__A1 _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5206__A2 _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4965__A1 _4206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8156__A1 _3208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7409__B _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7903__A1 _2961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9164__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5390__A1 _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7131__A2 _2291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5142__A1 _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5443__I _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5693__A2 _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6274__I _4418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7860_ _2369_ _2951_ _2987_ _2661_ _2988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_63_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8395__A1 _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6811_ _1987_ _2014_ _2022_ _2023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_91_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7791_ _2919_ _2920_ _2921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__6945__A2 _4176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6742_ _1954_ _1955_ _1956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_51_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8147__A1 _3175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6673_ _1900_ _1901_ _0083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5618__I _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8412_ _2196_ _2189_ _3428_ _3511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_34_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5624_ _0924_ _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8343_ _3293_ _3437_ _3443_ _3444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4803__S1 _4379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5555_ _0851_ _0626_ _0858_ _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5381__A1 _4155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7833__I _2961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8274_ _3376_ _3377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5486_ _0790_ _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7225_ _2369_ _2370_ _2371_ _0165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6449__I _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5133__A1 as2650.holding_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8870__A2 _3935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7156_ _2139_ _1921_ _2314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6107_ _1372_ _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8622__A2 _3345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7087_ _2197_ _2247_ _2250_ as2650.stack\[1\]\[5\] _2244_ _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_101_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5436__A2 _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6038_ _1303_ _0886_ _1304_ _1305_ _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__6484__I1 as2650.r123_2\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6184__I _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7189__A2 _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8386__A1 _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7989_ _2577_ _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_54_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__9187__CLK clknet_leaf_65_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8310__A1 _3082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8310__B2 _2645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6359__I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5124__B2 as2650.stack\[6\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8613__A2 _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5427__A2 _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6094__I _4194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8377__A1 _2482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6927__A2 _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7918__I _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8129__A1 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7352__A2 _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5340_ _0556_ _0557_ _0560_ _0567_ _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_115_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8301__A1 _2581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6269__I _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5271_ _0500_ _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7010_ _1118_ _1009_ _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8417__C _3154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6615__A1 as2650.r0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7958__A4 _3082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8961_ _3966_ _2129_ _4005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5969__A3 _4425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6091__A2 _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7912_ _1003_ _2525_ _3038_ _3001_ _3039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_71_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8892_ as2650.stack\[7\]\[11\] _3951_ _3954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_58_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7843_ _2969_ _2527_ _2970_ _2971_ _2972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_51_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6918__A2 _2114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_52_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7040__A1 _2201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7040__B2 as2650.stack\[4\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7774_ _1546_ _2903_ _2904_ _2905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4986_ as2650.holding_reg\[1\] _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6725_ _1716_ _1939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8135__A4 _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6656_ _1843_ _1884_ _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__8540__A1 _3076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5607_ _0909_ _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5354__A1 _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6587_ _0585_ _1721_ _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9375_ _0268_ clknet_leaf_75_wb_clk_i as2650.r123\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_69_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8326_ _2181_ _0919_ _3355_ _3427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_30_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5538_ _0517_ _0681_ _4546_ _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5106__A1 _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8257_ as2650.stack\[3\]\[1\] _4474_ _4473_ _3360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5469_ _0296_ _0740_ _0774_ _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5083__I _4312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7208_ _2357_ _2358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8188_ _3291_ _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7139_ _2300_ _2281_ _2283_ as2650.stack\[3\]\[4\] _2278_ _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_101_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_55_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_55_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_100_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output25_I net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9020__A2 _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7738__I _2868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6909__A2 _2019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7031__A1 _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6385__A3 _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5593__A1 _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5258__I _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9202__CLK clknet_leaf_47_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5721__I _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8598__A1 _3394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8598__B2 _3471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9352__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5877__B _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9011__A2 _4048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4840_ _4190_ _4421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9068__C _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7573__A2 _2707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8770__A1 _3842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4771_ _4304_ _4351_ _4352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_53_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6510_ as2650.r123\[0\]\[2\] as2650.r123_2\[0\]\[2\] as2650.psl\[4\] _1744_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7490_ _2178_ _2580_ _2626_ _2627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8522__A1 _3210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7325__A2 _2456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6441_ _0876_ _1682_ _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_70_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7383__I _2520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9160_ _0053_ clknet_leaf_58_wb_clk_i as2650.stack\[4\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5887__A2 _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6372_ _1520_ _1537_ _1628_ _1629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__9078__A2 _4105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8111_ _3164_ _3221_ _3067_ _3222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_138_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5323_ _4477_ _0629_ _0630_ _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_9091_ _4121_ _4122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8042_ _2440_ _2461_ _3155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6836__A1 _2021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5254_ _4338_ _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5185_ as2650.r123\[1\]\[4\] as2650.r123\[0\]\[4\] as2650.r123_2\[1\]\[4\] as2650.r123_2\[0\]\[4\]
+ _4196_ _0493_ _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__4942__S0 _4139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8053__A3 _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7986__C _2578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8944_ _3988_ _3993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4691__B _4271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8875_ _0938_ _3925_ _3942_ _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6462__I _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7826_ _2880_ _2952_ _2744_ _2955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7564__A2 _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8761__A1 _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7757_ _2485_ _2888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_36_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4969_ _4501_ _4540_ _4548_ _4549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_138_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6708_ as2650.stack\[0\]\[9\] _1927_ _1928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_137_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7688_ _2775_ _2797_ _2820_ _2821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5327__A1 _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9225__CLK clknet_leaf_55_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6639_ _1852_ _1854_ _1868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_137_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5878__A2 _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9358_ _0251_ clknet_leaf_59_wb_clk_i as2650.stack\[7\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__9069__A2 _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8309_ _0376_ _2533_ _1508_ _3410_ _3411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_133_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8816__A2 _3856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9289_ _0182_ clknet_leaf_28_wb_clk_i net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6827__A1 _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8292__A3 _3155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7252__A1 _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6055__A2 _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5566__A1 _4255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8504__A1 _3103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7307__A2 _4430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9335__D _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4620__I _4200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5869__A2 _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7931__I _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8807__A2 _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5652__S _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6975__C _2173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7491__A1 _2609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5451__I _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8762__I _4434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6990_ _2191_ _2164_ _2168_ as2650.stack\[2\]\[4\] _2142_ _2192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_66_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5941_ _0840_ _1165_ _1215_ _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_59_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7378__I _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5872_ _4527_ _1101_ _1150_ _1110_ _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_8660_ _4419_ _1046_ _4395_ _3749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_94_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7546__A2 _2580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8743__A1 _3827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7611_ _2704_ _2742_ _2743_ _2744_ _2745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_107_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4823_ _4364_ _4377_ _4403_ _4404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8591_ _2995_ _3621_ _3683_ _3592_ _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__9248__CLK clknet_leaf_63_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8711__B _3798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7542_ _2661_ _2677_ _2650_ _2479_ _2340_ _2678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_119_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4754_ _4332_ _4334_ _4309_ _4335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8430__C _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7473_ net29 _2417_ _2610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4685_ _4264_ _4265_ _4266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5626__I _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9212_ _0105_ clknet_leaf_75_wb_clk_i as2650.r123_2\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6424_ _1668_ _1660_ _1669_ _0066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9143_ _0036_ clknet_leaf_67_wb_clk_i as2650.r123_2\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6355_ _1253_ _1612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5306_ _0613_ _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_9074_ _4105_ _4108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6286_ _1335_ _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6285__A2 _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5237_ _0461_ _0371_ _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8025_ _3141_ _0637_ _3130_ _3142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5361__I _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5168_ _0354_ _4505_ _0369_ _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_84_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6037__A2 _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5099_ _0407_ _0310_ _0408_ _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8982__A1 _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8927_ _3978_ _3979_ _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5796__A1 _4406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6192__I _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8858_ _0848_ _3925_ _3930_ _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7537__A2 _2672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8734__A1 _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7809_ _2924_ _2933_ _2938_ _2939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XPHY_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8789_ _0711_ _3856_ _3245_ _3873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5720__A1 _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5720__B2 as2650.r123_2\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6367__I _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6276__A2 _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5271__I _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7225__A1 _2369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4615__I _4138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8025__I0 _3141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5539__A1 _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6200__A2 _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5446__I _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4762__A2 _4311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7700__A2 _2809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7661__I _2793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6140_ _1399_ _0681_ _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7464__A1 as2650.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6277__I _4227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6071_ _1322_ _1086_ _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5022_ as2650.stack\[0\]\[9\] _4465_ _0324_ as2650.stack\[1\]\[9\] _0333_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_79_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7216__A1 _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6973_ _2174_ _2177_ _0107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8712_ _3199_ _4535_ _3789_ _3799_ _3800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5924_ _0749_ _1057_ _1145_ _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7519__A2 _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8716__A1 _3703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8643_ _3430_ _3730_ _3732_ _2482_ _3733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_110_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5855_ _0389_ _1097_ _1134_ _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6578__I0 as2650.r123\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4806_ _4386_ _4387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8574_ _0996_ _3666_ _3667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_124_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5786_ _1067_ _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7525_ _2336_ _2479_ _2661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4737_ _4317_ _4311_ _4318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_120_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7456_ _4511_ _4512_ _4528_ _2593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4668_ as2650.ins_reg\[4\] _4249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_6407_ _1655_ _1656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7387_ _2524_ _2525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4599_ as2650.ins_reg\[2\] _4180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9126_ _0019_ clknet_leaf_59_wb_clk_i as2650.stack\[6\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6338_ as2650.psl\[5\] _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_1_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7455__A1 _4503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7455__B2 _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6269_ _1280_ _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9057_ _3851_ _1100_ _4092_ _4093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8008_ _1699_ _1295_ _3128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7207__A1 _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7758__A2 _2883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8955__A1 _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5233__A3 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6430__A2 _1661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8707__A1 _4458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6194__A1 _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5941__A1 _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4744__A2 _4324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7694__A1 _2825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7481__I _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7414__C _2551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6249__A2 _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7446__A1 _2581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7749__A2 _2878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4680__A1 _4250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5640_ as2650.pc\[5\] _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__7921__A2 _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5571_ _0874_ _4193_ _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7310_ _0469_ _1261_ _4425_ _2449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_116_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8290_ _1267_ _3057_ _3155_ _1288_ _3392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_117_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7241_ _2382_ _2383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7172_ _2298_ _2322_ _2327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7437__A1 _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6123_ _0464_ _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7988__A2 _3107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6054_ _1326_ _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5005_ _4332_ _4386_ _4324_ _0315_ _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_113_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4671__A1 as2650.cycle\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8155__C _3207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6956_ _0969_ _2161_ _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5907_ _0505_ _1066_ _1183_ _1076_ _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6887_ _2093_ _2096_ _2097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_22_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8165__A2 _3074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8626_ _2926_ _3706_ _3716_ _3598_ _3717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6176__A1 _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5838_ _1089_ _1118_ _4444_ _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__7373__B1 _2502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7912__A2 _2525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8557_ _1709_ _2976_ _3650_ _3651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5923__A1 _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5086__I _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5769_ _1038_ _1039_ _1041_ _1050_ _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_124_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7508_ _1579_ _2644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8488_ as2650.stack\[7\]\[7\] _3366_ _3361_ as2650.stack\[4\]\[7\] as2650.stack\[5\]\[7\]
+ _3362_ _3585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8397__I _3495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7439_ _1390_ _2577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5814__I _4233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4858__C _4438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7428__A1 _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9109_ _0002_ clknet_leaf_68_wb_clk_i as2650.r123\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5035__B _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4874__B _4454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6651__A2 _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5689__C _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8928__A1 _3976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9050__B1 _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8860__I _3928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5057__I3 as2650.r123_2\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7476__I _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4965__A2 _4543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8156__A2 _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6167__A1 as2650.stack\[4\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9309__CLK clknet_leaf_16_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7144__C _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7419__A1 _4529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8092__A1 _3136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6642__A2 _1849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8919__A1 _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5996__A4 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6810_ _1989_ _2013_ _2022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_42_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7790_ net36 _2885_ _2920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6741_ _0672_ _1732_ _1878_ _1955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_32_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4956__A2 _4535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8147__A2 _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7386__I _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6158__A1 _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6672_ _1223_ _1717_ _1901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8411_ _2736_ _2756_ _3504_ _3509_ _3510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_104_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5905__A1 _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5623_ _0535_ _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8342_ _2854_ _3425_ _3442_ _3058_ _3443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5554_ _0857_ _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5381__A2 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4959__B _4537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7658__A1 _2778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8273_ _3055_ _3284_ _3285_ _3286_ _3376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_5485_ _0789_ _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8010__I _3119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7224_ _1556_ _2359_ _2371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5133__A2 _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7155_ _2312_ _2313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8083__A1 _2383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6106_ _4441_ _1376_ _1378_ _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7086_ _2186_ _2245_ _2263_ _0134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6465__I _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6037_ _4254_ _0878_ _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4644__A1 _4159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7189__A3 _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8680__I _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6397__A1 _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7988_ _4243_ _3107_ _3111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6939_ _2144_ _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4713__I _4285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7897__A1 _2998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8609_ _3210_ _3686_ _3700_ _3701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7649__A1 _2777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5544__I _4295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6321__A1 _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8613__A3 _3663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7821__A1 _2899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5212__C _4247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8377__A2 _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9131__CLK clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4938__A2 _4517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8129__A2 _2658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7888__A1 as2650.pc\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9281__CLK clknet_leaf_26_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8031__S _3130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8301__A2 _4380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5270_ _0577_ _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_9_wb_clk_i_I clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5115__A2 _4452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8960_ _0775_ _3986_ _3989_ as2650.r123\[2\]\[6\] _4004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_56_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4626__A1 _4163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7911_ _3035_ _2495_ _3036_ _3037_ _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_110_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8891_ _1666_ _3948_ _3953_ _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_37_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7842_ net53 _2531_ _2535_ _2366_ _2854_ _2971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__6379__A1 _1611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7773_ _2884_ _2618_ _2500_ _2904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4985_ _0295_ _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6724_ _1937_ _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7879__A1 _2982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6655_ _1880_ _1881_ _1883_ _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_5606_ as2650.pc\[1\] _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5792__C _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9374_ _0267_ clknet_leaf_77_wb_clk_i as2650.r123\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5354__A2 _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6586_ _1758_ _1805_ _1816_ _1777_ _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_121_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8325_ _2387_ _3426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5537_ _0839_ _0841_ _4364_ _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5364__I as2650.r0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8256_ _3338_ _3343_ _3352_ _3358_ _3359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6303__A1 _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5468_ _0285_ _0749_ _0773_ _0295_ _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_82_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7207_ _1569_ _2339_ _2344_ _2356_ _2357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_78_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8187_ _3290_ _3291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5399_ as2650.stack\[0\]\[13\] _4481_ _0324_ as2650.stack\[1\]\[13\] _0706_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_120_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8056__A1 _1612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7138_ _2190_ _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7803__A1 _2514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4708__I _4288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7069_ _2147_ _2247_ _2250_ as2650.stack\[1\]\[0\] _2244_ _2251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_74_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4617__A1 _4197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7567__B1 _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7031__A2 _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output18_I net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_24_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_24_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5593__A2 _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8531__A2 _3610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5345__A2 _4191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8295__A1 _3395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8518__C _2928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8047__A1 _3158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4618__I _4198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4608__A1 _4161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5449__I net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5033__A1 _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4770_ _4348_ _4350_ _4351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8522__A2 _3596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7325__A3 _2463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6440_ _4223_ _1681_ _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5184__I _4379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6371_ _1480_ _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8110_ _2151_ _3221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5322_ as2650.stack\[7\]\[12\] _4479_ _4461_ as2650.stack\[6\]\[12\] _0630_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8286__A1 _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9090_ _4065_ _4120_ _4121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_114_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8709__B _1480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8041_ _2149_ _3154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8495__I _2577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5253_ _0560_ _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8428__C _3526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5184_ _4379_ _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_64_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4942__S1 _4379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7261__A2 _2401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6064__A3 _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8943_ _3986_ _3992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8444__B _3181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8874_ _2302_ _3927_ _3929_ as2650.stack\[7\]\[5\] _3924_ _3942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__8210__A1 _2335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7825_ _2336_ _2612_ _2952_ _2953_ _2954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_51_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8761__A2 _3772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7756_ _2480_ _2886_ _2887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4968_ _4542_ _4547_ _4548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6707_ _1922_ _1927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7687_ _2751_ _2813_ _2819_ _2820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4899_ as2650.stack\[7\]\[8\] _4479_ _4461_ as2650.stack\[6\]\[8\] _4480_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8513__A2 _3566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6638_ _1836_ _1857_ _1866_ _1867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_137_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9357_ _0250_ clknet_leaf_60_wb_clk_i as2650.stack\[7\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6569_ _1799_ _1789_ _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8308_ _2365_ _2754_ _3410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_9288_ _0181_ clknet_leaf_27_wb_clk_i net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8239_ _2777_ _3340_ _3341_ _3089_ _3342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_133_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8029__A1 _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7252__A2 _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6460__B1 _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8201__A1 _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6763__A1 _1949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5566__A2 _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8504__A2 _3598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7307__A3 _4432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4901__I _4481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7433__B _2570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7491__A2 _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8440__A1 _2800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5940_ _0516_ _1164_ _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5871_ _0566_ _1103_ _1127_ _1149_ _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_61_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7610_ _1341_ _2744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8743__A2 _3773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4822_ _4378_ _4388_ _4402_ _4222_ _4403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_8590_ _3292_ _3665_ _3682_ _3331_ _3683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8711__C _3765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9095__B net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7541_ _2670_ _2676_ _2677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4753_ _4333_ _4334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7394__I _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4811__I _4391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7472_ net30 _2609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4684_ as2650.addr_buff\[5\] _4265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_9211_ _0104_ clknet_leaf_76_wb_clk_i as2650.r123_2\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6423_ as2650.stack\[2\]\[11\] _1664_ _1669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_128_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9142_ _0035_ clknet_leaf_67_wb_clk_i as2650.r123_2\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6354_ as2650.psl\[7\] _1611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5305_ _0610_ _0503_ _0572_ _0611_ _0612_ _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_9073_ _1089_ _4106_ _4107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6285_ _1522_ _1542_ _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8024_ _1290_ _3140_ _3141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5236_ _4325_ _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5167_ _0475_ _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_5_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5798__B _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5098_ _0402_ _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7569__I _2703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6473__I _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8982__A2 _3236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8926_ _0703_ _3969_ _3979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8857_ _2146_ _3927_ _3929_ as2650.stack\[7\]\[0\] _3924_ _3930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XPHY_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7808_ _2377_ _2936_ _2937_ _2938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8788_ _3861_ _3871_ _3872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7739_ _2866_ _2867_ _2869_ _2870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_123_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9342__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5720__A2 _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7473__A2 _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8670__A1 _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7225__A2 _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8422__B2 _4453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8084__B _3195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6383__I _1638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8973__A2 _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6316__C _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8025__I1 _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8812__B _1629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6736__A1 _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5539__A2 _4547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8103__I _3045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7147__C _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7464__A2 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6070_ _1339_ _1342_ _1323_ _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8661__A1 _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8661__B2 _3265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input9_I io_in[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5475__B2 _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5021_ as2650.stack\[2\]\[9\] _4460_ _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8413__A1 _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7216__A2 _2358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7389__I _2526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5227__A1 _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9215__CLK clknet_leaf_41_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6293__I _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4806__I _4386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6972_ _0908_ _2176_ _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6975__A1 _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6226__C _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8711_ _3790_ _0400_ _3798_ _3765_ _3799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_111_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5923_ _0771_ _1097_ _1134_ _1198_ _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_94_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8642_ _4264_ _2410_ _2494_ _3726_ _3731_ as2650.pc\[14\] _3732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_34_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6727__A1 _1939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5854_ _1133_ _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_80_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9365__CLK clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6578__I1 as2650.r123_2\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4805_ _4381_ _4385_ _4386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_8573_ _0989_ _3648_ _3666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5785_ _4228_ _1042_ _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7524_ _2638_ _2659_ _2660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4736_ as2650.psl\[3\] _4316_ _4317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5950__A2 _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7455_ _4503_ _0350_ _0356_ _0386_ _0387_ _2592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
X_4667_ _4149_ _4248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6406_ _1654_ _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7386_ _2523_ _2524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4598_ _4178_ _4179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_115_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6468__I _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9125_ _0018_ clknet_leaf_57_wb_clk_i as2650.stack\[6\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6337_ _1585_ _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5372__I _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7455__A2 _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9056_ _1627_ _0818_ _3115_ _4091_ _1628_ _4092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_6268_ _0758_ _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_103_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5466__A1 _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8007_ _0361_ _3126_ _3127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5219_ as2650.stack\[3\]\[11\] _4450_ _4469_ as2650.stack\[1\]\[11\] _0528_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_131_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6199_ _0394_ _1452_ _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8404__A1 _3221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7299__I _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4716__I _4280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5769__A2 _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8909_ _3961_ _3966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8707__A2 _3793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8183__A3 _3285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7391__A1 _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6194__A2 _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5547__I _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5941__A2 _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5991__B _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7143__A1 _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7694__A2 _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8891__A1 _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6351__C1 _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6378__I _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7446__A2 _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8643__B2 _2482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5457__A1 _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9238__CLK clknet_leaf_39_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5209__A1 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4680__A2 _4151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9388__CLK clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6709__A1 _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7921__A3 _3046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5570_ _4184_ _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7134__A1 _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7134__B2 as2650.stack\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7240_ _1479_ _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7171_ _2296_ _2318_ _2319_ as2650.stack\[0\]\[3\] _2320_ _2326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_131_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6122_ _1373_ _1388_ _1389_ _1392_ _0041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7437__A2 _2522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_71_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6053_ _0883_ _1325_ _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5004_ _0297_ _0314_ _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4671__A2 as2650.cycle\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6955_ _2149_ _0875_ _2159_ _0897_ _2160_ _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_54_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6751__I _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5906_ _0718_ _1068_ _1069_ _1182_ _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6886_ _2094_ _2095_ _2096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8625_ _2372_ _3669_ _3500_ _2382_ _3716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5837_ _0969_ _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6176__A2 _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8556_ _0990_ _1544_ _3650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5768_ _1042_ _1046_ _1049_ _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_72_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7507_ net31 _2643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4719_ _4286_ _4300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8678__I _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8487_ as2650.stack\[0\]\[7\] _1905_ _1657_ as2650.stack\[1\]\[7\] _0525_ _3584_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5699_ _0992_ _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7438_ _2530_ _2520_ _2576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7676__A2 _2741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8873__A1 _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6333__C1 _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_49_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_104_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7369_ _2507_ _2508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9108_ _0001_ clknet_leaf_68_wb_clk_i as2650.r123\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8625__A1 _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5439__A1 _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9039_ _3088_ _0570_ _4076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8928__A2 _1859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9050__A1 _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9050__B2 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8362__B _1685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7757__I _2485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4965__A3 _4544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6167__A2 _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5277__I as2650.r0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8864__A1 _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5678__A1 as2650.r123\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8616__A1 _3035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7419__A2 _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8092__A2 _3061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5850__A1 _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8919__A2 _3959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8395__A3 _3423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7667__I _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5602__A1 _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6740_ _1847_ _1953_ _1954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_51_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9087__C _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6671_ as2650.r123_2\[1\]\[7\] _1729_ _1899_ _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_108_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8410_ _2509_ _3508_ _3509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5622_ _0923_ _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9390_ _0283_ clknet_leaf_5_wb_clk_i as2650.psu\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5905__A2 _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8341_ _3181_ _3440_ _3441_ _2925_ _3442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5553_ _0856_ _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7658__A2 _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8272_ _3333_ _3335_ _3372_ _3374_ _3375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_144_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5484_ _0788_ _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7223_ _2357_ _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6866__B1 _2076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8607__A1 _3458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7154_ _0851_ _1921_ _2162_ _2312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_141_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4892__A2 _4450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6105_ _1377_ _1100_ _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8083__A2 _3061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7085_ _2191_ _2247_ _2250_ as2650.stack\[1\]\[4\] _2244_ _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__5650__I _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6036_ _0888_ _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7830__A2 _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4644__A2 _4179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9032__A1 _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7594__A1 _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7987_ _4264_ _2824_ _3110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6397__A2 _1643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6938_ _0862_ _2144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6149__A2 _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7346__A1 _2484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6869_ _2078_ _2079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_50_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8608_ _0632_ _1499_ _3699_ _3700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7897__A2 _2876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8539_ _2526_ _3623_ _3633_ _1234_ _3634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_109_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7649__A2 _2780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8846__A1 _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4580__A1 _4157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5109__C2 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6321__A2 _4314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4883__A2 _4463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8074__A2 _3186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5560__I _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6085__A1 _4551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7821__A2 _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5832__A1 _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9023__A1 _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7487__I _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4904__I _4445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4874__A2 _4452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6076__A1 as2650.cycle\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4626__A2 _4165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7910_ net52 _2504_ _2507_ _3020_ _1268_ _3037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__9014__A1 _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8890_ as2650.stack\[7\]\[10\] _3951_ _3953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7025__B1 _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7841_ _2540_ _2947_ _2970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7397__I _2534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6379__A2 _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7772_ _2890_ _2902_ _2903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4984_ _0294_ _4261_ _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_23_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6723_ _1934_ _1936_ _1261_ _1937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7879__A2 _2644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6654_ as2650.r0\[0\] _1882_ _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6000__A1 _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8540__A3 _3634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5605_ _0337_ _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9373_ _0266_ clknet_leaf_74_wb_clk_i as2650.r123\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6585_ _1759_ _1746_ _1783_ _1757_ _1816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_121_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8324_ _3424_ _3425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5536_ _4515_ _0840_ _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8255_ _3354_ _3335_ _3357_ _1289_ _3358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_106_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5467_ _4354_ _0768_ _0772_ _0700_ _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_65_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7500__A1 _2181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7206_ _2351_ _2355_ _1701_ _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_114_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8186_ _1358_ _3290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5398_ as2650.stack\[6\]\[13\] _4461_ _0329_ _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7137_ _2297_ _2299_ _0149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8056__A2 _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6476__I _1712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7068_ _2249_ _2250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4617__A2 _4135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9005__A1 _2635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8691__I _4394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6019_ _4443_ _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7567__A1 _2190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6144__C _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8516__B1 _3611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_64_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_64_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_52_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8819__A1 _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7703__C _2476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5290__I _4396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6058__A1 _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5805__A1 _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4608__A2 _4171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7558__A1 _2687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4634__I _4181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6230__A1 _1486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5584__A3 _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6070__B _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5465__I _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7730__A1 _2751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6370_ _1519_ _1627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_127_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5321_ as2650.stack\[4\]\[12\] _4482_ _0626_ as2650.stack\[5\]\[12\] _0629_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_115_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8040_ _1685_ _3153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5252_ _4488_ _0504_ _0559_ _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6296__I _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4809__I net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5183_ _0364_ _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6064__A4 _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8942_ _4414_ _3987_ _3990_ _3991_ _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_83_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8873_ _0932_ _3925_ _3941_ _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_97_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7824_ _2871_ _2869_ _2564_ _2953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7755_ _2884_ _2885_ _2886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_36_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4967_ _4546_ _4547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6706_ _1653_ _1924_ _1926_ _0091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7686_ _2613_ _2780_ _2817_ _2818_ _2819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_32_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4898_ _4478_ _4479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_123_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6637_ _1837_ _1856_ _1866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5375__I net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7721__A1 net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6568_ _1779_ _1787_ _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_9356_ _0249_ clknet_leaf_59_wb_clk_i as2650.stack\[7\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8307_ _1336_ _2620_ _3408_ _3409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5519_ _0599_ _0744_ _0717_ _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_9287_ _0180_ clknet_leaf_27_wb_clk_i net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6499_ _4541_ _1733_ _1724_ _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_8238_ _4530_ _2503_ _3341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9121__CLK clknet_leaf_39_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4719__I _4286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8029__A2 _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8169_ _0867_ _0879_ _1682_ _2346_ _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_47_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6139__C _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7788__A1 _2476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7788__B2 _2554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7252__A3 _2393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8354__C _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6460__A1 _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6460__B2 _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6212__A1 _4543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7960__A1 _3080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8504__A3 _3353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7307__A4 _1470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5285__I _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7005__I _2203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7779__A1 _2884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8440__A2 _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5888__C _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8264__C _4476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6451__A1 _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5870_ _0512_ _1146_ _1148_ _1102_ _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_34_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6203__A1 _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4821_ _4389_ _4401_ _4402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7540_ _1594_ _2473_ _2675_ _2564_ _2676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4752_ _4304_ _4333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_109_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7471_ _2602_ _2605_ _2607_ _2608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4683_ as2650.addr_buff\[6\] _4264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5195__I _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7703__A1 _2704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9210_ _0103_ clknet_leaf_77_wb_clk_i as2650.r123_2\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6422_ _0999_ _1668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9141_ _0034_ clknet_leaf_67_wb_clk_i as2650.r123_2\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6353_ _1261_ _1527_ _1603_ _1609_ _1610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_66_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5304_ _0348_ _0574_ _0575_ _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_143_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9072_ _2373_ _3144_ _4105_ _4106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6284_ _1045_ _1534_ _1536_ _1539_ _1541_ _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__9294__CLK clknet_leaf_25_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8023_ _2736_ _3103_ _3140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5235_ as2650.holding_reg\[4\] _0542_ _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_64_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6690__A1 _1668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5166_ _0446_ _0474_ _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5097_ _0303_ _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_83_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8925_ as2650.r123\[1\]\[5\] _3967_ _3977_ _3978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_71_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8856_ _3928_ _3929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8195__A1 _2899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7807_ _2919_ _2644_ _2852_ _2937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7585__I _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7942__A1 _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5999_ _1243_ _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8787_ _0690_ _2633_ _3870_ _2630_ _3871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7738_ _2868_ _2869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8498__A2 _3561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7669_ _2799_ _2734_ _2801_ _2802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_138_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7534__B _2662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5181__A1 _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9339_ _0232_ clknet_leaf_51_wb_clk_i as2650.stack\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8349__C _4475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8670__A2 _4361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8422__A2 _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6433__A1 _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7709__B _2818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7495__I _2443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6736__A2 _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7428__C _2565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9167__CLK clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_61_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8661__A2 _3748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6672__A1 _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5020_ as2650.stack\[3\]\[9\] _4452_ _4454_ _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8275__B _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8949__B1 _3993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6424__A1 _1668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6971_ _2175_ _2140_ _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_65_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6975__A2 _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8710_ _3791_ _3796_ _3797_ _3798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5922_ _1099_ _1196_ _1197_ _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_81_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8177__A1 _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8641_ _3081_ _3731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5853_ _4552_ _1037_ _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7924__A1 _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6727__A2 _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4804_ _4383_ _4140_ _4286_ _4384_ _4385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__4738__A1 _4315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8572_ _3664_ _3665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5935__B1 _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5784_ _1065_ _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7523_ _2639_ _2606_ _2659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4735_ as2650.carry _4316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_30_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7454_ _1699_ _2553_ _2467_ _2590_ _2591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4666_ _4233_ _4206_ _4242_ _4246_ _4247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_31_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6405_ _4456_ as2650.psu\[1\] _1654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5163__A1 _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5163__B2 _4225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7385_ _1498_ _4418_ _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4597_ _4177_ _4178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_9124_ _0017_ clknet_leaf_57_wb_clk_i as2650.stack\[6\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6336_ _1523_ _1578_ _1592_ _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8101__A1 _3209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9055_ _4072_ _3113_ _1519_ _4091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_130_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6267_ as2650.psl\[6\] _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5466__A2 _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5218_ _0426_ _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_8006_ _1289_ _3126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6198_ _1454_ _1455_ _0789_ _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_130_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8404__A2 _3499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5149_ _4518_ _0457_ _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5769__A3 _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8908_ _4414_ _3959_ _3965_ _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4977__A1 _4305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8168__A1 _3262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8839_ _2298_ _3912_ _3917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7915__A1 _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6718__A2 _1923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7915__B2 _2940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4729__A1 _4256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7391__A2 _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7930__A4 _3055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5991__C _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8340__A1 _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8891__A2 _3948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6351__B1 _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5563__I _4214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6351__C2 _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7446__A3 _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6654__A1 as2650.r0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8095__B _3189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4907__I _4191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5209__A2 _4526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4680__A3 _4260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6957__A2 _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4968__A1 _4542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8159__A1 _3263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7906__A1 _2607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7921__A4 _2433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8331__A1 _2182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7134__A2 _2286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6893__A1 _1174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7170_ _2324_ _2325_ _0156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6121_ _1391_ _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6645__A1 _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7842__B1 _2535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6052_ _4174_ _4207_ _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5422__B _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5003_ _4331_ _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8398__A1 _3393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9332__CLK clknet_leaf_80_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7070__A1 _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6954_ _0898_ _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5905_ _0690_ _1146_ _1181_ _1102_ _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_81_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5648__I _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6885_ _2028_ _2071_ _2095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8624_ _3093_ _3714_ _3715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5836_ _1090_ _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7373__A2 _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5384__A1 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8555_ _2969_ _3648_ _3649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5767_ _1047_ _1048_ _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7506_ _1614_ _2641_ _2642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_108_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4718_ _4298_ _4281_ _4299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_136_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8322__A1 as2650.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5698_ _0990_ _0980_ _0973_ as2650.r123_2\[0\]\[2\] _0991_ _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_8486_ as2650.stack\[3\]\[7\] _1920_ _1639_ as2650.stack\[2\]\[7\] _3583_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_7437_ _0912_ _2522_ _2574_ _2575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4649_ _4229_ _4230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6333__B1 _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6333__C2 _4392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7368_ _2506_ _2507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9107_ _0000_ clknet_leaf_66_wb_clk_i as2650.r123\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6319_ _1575_ _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8625__A2 _3669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7299_ _0869_ _2438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8627__C _2856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9038_ _3851_ _4074_ _3868_ _4075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_18_wb_clk_i clknet_3_3_0_wb_clk_i clknet_leaf_18_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_131_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8389__A1 _3481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__9050__A2 _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6942__I _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7061__A1 _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5558__I as2650.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9177__D _0070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8561__A1 _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5127__A1 _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9205__CLK clknet_leaf_74_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8864__A2 _3935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6875__A1 _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5678__A2 _4153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8616__A2 _3687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9355__CLK clknet_leaf_60_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7441__C _2578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8272__C _3374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5602__A2 _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6670_ _1795_ _1898_ _1899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_43_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8552__A1 _2952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5621_ _0918_ _0922_ _0915_ _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_143_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5366__A1 _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8340_ _1147_ _3157_ _3441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5552_ _0852_ _0855_ _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7616__C _2658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8304__A1 _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8271_ _3373_ _3374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5118__A1 as2650.stack\[2\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5483_ _4367_ _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8855__A2 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7222_ _2368_ _2369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6866__B2 _1980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7153_ _2310_ _2311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8607__A2 _3686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4975__C _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6618__A1 _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6104_ _1375_ _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7084_ _2261_ _2262_ _0133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8083__A3 _3192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6035_ _4263_ _1307_ _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7291__A1 _1939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5841__A2 _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7043__A1 _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7986_ _3107_ _3108_ _3109_ _2578_ _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7594__A2 _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8791__A1 _2565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6937_ _2142_ _2143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5378__I _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6868_ _2062_ _2065_ _2078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_74_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7346__A2 _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8543__A1 _3257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8543__B2 _2549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7807__B _2852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8607_ _3458_ _3686_ _3698_ _3699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9228__CLK clknet_leaf_40_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5819_ _4334_ _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_91_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7897__A3 _2878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6799_ _2003_ _2011_ _2012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8538_ _1275_ _3341_ _3632_ _3633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_109_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5109__A1 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5109__B2 _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8469_ _3564_ _3540_ _3565_ _3566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_68_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4580__A2 _4160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6002__I _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8638__B _3625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6321__A3 _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6609__A1 _4382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7282__A1 _4551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6085__A2 _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7821__A3 _2366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9023__A2 _4059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7768__I _2866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7034__A1 _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8782__A1 _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5596__A1 _4152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5288__I _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8534__A1 _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5348__A1 _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4920__I _4274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6340__C _1596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6848__A1 _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7452__B _2588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5520__A1 _4374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7171__C _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7273__A1 _2403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4706__S0 as2650.ins_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7025__A1 _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7840_ _2968_ _2969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_37_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8773__A1 _3837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5587__A1 _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7771_ _2785_ _2891_ _2893_ _2902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5198__I _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4983_ _4248_ _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6722_ _1038_ _1215_ _1133_ _1935_ _1936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_108_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7627__B _2728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5339__A1 _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6653_ as2650.r123\[0\]\[7\] as2650.r123_2\[0\]\[7\] _4144_ _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6000__A2 _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5604_ _0848_ _0861_ _0907_ _0008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_9372_ _0265_ clknet_leaf_76_wb_clk_i as2650.r123\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6584_ _4383_ _1781_ _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8323_ _0927_ _3423_ _3424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5535_ _4320_ _4334_ _4321_ _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8254_ _3355_ _3356_ _3354_ _3357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5466_ _0486_ _0771_ _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7500__A2 _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7205_ _1524_ _2353_ _2354_ _2355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5511__A1 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8185_ _3288_ _3289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5397_ as2650.stack\[7\]\[13\] _0326_ _4466_ as2650.stack\[4\]\[13\] as2650.stack\[5\]\[13\]
+ _4470_ _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__5661__I _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8177__C _3280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7136_ _2298_ _2291_ _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_87_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7264__A1 _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7067_ _2165_ _2248_ _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6018_ _1291_ _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9005__A2 _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7567__A2 _2686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8764__A1 _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7969_ _3093_ _2155_ _2508_ _3094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8516__A1 _3598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8516__B2 _3070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5502__A1 _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7255__A1 _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8882__I _3946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5805__A2 _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7498__I _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7007__A1 _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7558__A2 _2532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8755__A1 _2477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5569__A1 _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6230__A2 _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8507__A1 _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4792__A2 _4372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5741__A1 _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5320_ _0623_ _0625_ _0627_ _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_142_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5251_ _0549_ _4421_ _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5481__I as2650.r123\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5182_ _0490_ _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8994__A1 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8941_ _3966_ _1979_ _3991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4825__I _4405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8872_ _2300_ _3927_ _3929_ as2650.stack\[7\]\[4\] _3924_ _3941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__8746__A1 _3810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7823_ _2866_ as2650.addr_buff\[1\] _2952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7754_ _2838_ _2839_ _2885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4966_ _4545_ _4546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8460__C _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6705_ as2650.stack\[0\]\[8\] _1925_ _1926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7685_ _2485_ _2818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5980__A1 as2650.psl\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4897_ _4450_ _4478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_36_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4560__I _4140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6636_ _1827_ _1863_ _1864_ _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7721__A2 _2644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9355_ _0248_ clknet_leaf_60_wb_clk_i as2650.stack\[7\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6567_ _1774_ _1796_ _1797_ _1798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_121_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8306_ _0919_ _1708_ _3408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5518_ _0611_ _0822_ _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9286_ _0179_ clknet_leaf_27_wb_clk_i net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6498_ _1732_ _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7485__A1 _2609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8237_ _4530_ _4380_ _3339_ _3340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_5449_ net2 _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5391__I _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8168_ _3262_ _3208_ _3229_ _3272_ _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_120_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7237__A1 _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7119_ _2138_ _2279_ _2284_ _0146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8099_ _3046_ _3210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8985__A1 _3415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_12_wb_clk_i_I clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5799__A1 _4353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4735__I as2650.carry vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6460__A2 _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output23_I net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6212__A2 _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5971__A1 _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7712__A2 _2816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_51_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8673__B1 _3183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7228__A1 _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8976__A1 _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6451__A2 _1692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8728__A1 _3769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8728__B2 _4435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8561__B _3654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5006__A3 _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4820_ _4392_ _4397_ _4400_ _4401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5962__A1 _4426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4751_ _4331_ _4332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8200__I0 _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7470_ _1338_ _2607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4682_ _4235_ _4236_ _4240_ _4263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__8900__A1 _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6421_ _1666_ _1660_ _1667_ _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_70_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6911__B1 _1942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9140_ _0033_ clknet_leaf_46_wb_clk_i as2650.r123_2\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7624__C _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6352_ _1606_ _1607_ _1608_ _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_127_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7467__A1 _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5303_ _4348_ _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9071_ _1270_ _1274_ _4103_ _4104_ _4105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_6283_ _1540_ _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6100__I _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8022_ _3139_ _0194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5234_ _0541_ _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_142_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7219__A1 _2366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6690__A2 _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5165_ _0397_ _0442_ _0455_ _0472_ _0473_ _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_68_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8967__A1 _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5096_ _0402_ _0405_ _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_68_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4555__I _4135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8924_ _3976_ _1823_ _3977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_44_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8027__I _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8719__A1 _3804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8855_ _2148_ _0624_ _0901_ _3928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_52_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8195__A2 _2755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7806_ _2912_ _2935_ _2936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_129_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8786_ _1292_ _3766_ _3869_ _3870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5998_ _1271_ _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_40_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7737_ _0836_ _0827_ _4245_ _2868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5953__A1 _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4949_ _4528_ _4529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7668_ _2800_ _0667_ _2801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_32_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8697__I _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6619_ _1844_ _1848_ _1849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_123_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7599_ _2694_ _0613_ _2733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9338_ _0231_ clknet_leaf_39_wb_clk_i as2650.stack\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5181__A2 _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9269_ _0162_ clknet_leaf_14_wb_clk_i as2650.addr_buff\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8365__C _2927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8958__A1 _3995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7630__A1 _2757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6433__A2 _1661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6680__I _1907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6197__A1 _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7697__A1 _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7449__A1 _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7016__I _2213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6672__A2 _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8949__A1 _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6970_ _0858_ _2175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_4_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5921_ _0751_ _1063_ _1061_ _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8177__A2 _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8640_ as2650.pc\[14\] _3729_ _3730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_80_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5852_ _0360_ _1099_ _1131_ _1061_ _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6188__A1 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9111__CLK clknet_leaf_68_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7924__A2 _2412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4803_ as2650.r123\[1\]\[1\] as2650.r123\[0\]\[1\] as2650.r123_2\[1\]\[1\] as2650.r123_2\[0\]\[1\]
+ _4139_ _4379_ _4384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_8571_ _0996_ _3663_ _3664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5783_ _4220_ _1042_ _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5935__B2 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7522_ _2340_ _2658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4734_ _4312_ _4314_ _4315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_72_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7453_ _2584_ _2587_ _2589_ _2590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4665_ _4245_ _4246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__9261__CLK clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6404_ _0975_ _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7384_ _2517_ _2522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5163__A2 _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4596_ as2650.ins_reg\[7\] _4177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9123_ _0016_ clknet_leaf_58_wb_clk_i as2650.stack\[6\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6335_ as2650.psu\[7\] _1579_ _1582_ as2650.psu\[4\] _1591_ _1592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_131_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8101__A2 _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9054_ _0821_ _1431_ _1518_ _4090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6266_ _1288_ _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_103_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8005_ _3125_ _0191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7860__A1 _2369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5217_ _0525_ _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_135_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6197_ _0751_ _0669_ _0500_ _0492_ _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_69_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5148_ _0359_ _4142_ _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5079_ _0385_ _0388_ _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_44_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8907_ _3962_ _1724_ _3964_ as2650.r123\[1\]\[0\] _3965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_25_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4977__A2 _4306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8168__A2 _3208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8838_ _2296_ _3908_ _3909_ as2650.stack\[6\]\[3\] _3910_ _3916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__7376__B1 _2512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7915__A2 _2522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5926__A1 _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4729__A2 _4304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8769_ _0603_ _2633_ _3853_ _3854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7679__A1 _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5844__I _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8340__A2 _3157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6351__A1 _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6351__B2 _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8376__B _3475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7851__A1 _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6654__A2 _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6675__I _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7851__B2 _2940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7603__A1 _2736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9134__CLK clknet_leaf_56_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6957__A3 _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4968__A2 _4547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8159__A2 _3074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9000__B _4026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7906__A2 _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5917__A1 _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9284__CLK clknet_leaf_26_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8331__A2 _1617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6893__A2 _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6120_ _1390_ _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7902__C _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7842__A1 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6051_ _0889_ _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7842__B2 _2366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5002_ _4277_ _4329_ _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6953_ _2152_ _2158_ _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4959__A2 _4527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5904_ _1180_ _1146_ _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6884_ _2057_ _2070_ _2094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8623_ _3710_ _3711_ _3713_ _3714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5835_ _1094_ _1114_ _1115_ _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5908__A1 _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8570__A2 _3644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8554_ _3620_ _3597_ _3648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5766_ _4195_ _1042_ _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5384__A2 _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7505_ _2638_ _2640_ _2641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4717_ _4297_ _4298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8485_ _2492_ _3574_ _3581_ _3001_ _3582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5697_ _0347_ _0981_ _0982_ _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8322__A2 _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8040__I _1685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7436_ _2552_ _2572_ _2573_ _2574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4648_ _4212_ _4228_ _4229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6333__A1 as2650.psu\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6333__B2 net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7367_ _0881_ _2154_ _2506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_122_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4579_ _4159_ _4160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9106_ _4132_ _4134_ _1302_ _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8086__A1 _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6318_ _1374_ _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_46_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7298_ _1497_ _4543_ _2437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9037_ _1627_ _0566_ _3141_ _4073_ _4074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_77_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6249_ _1464_ _0883_ _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_104_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4647__A1 _4223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8389__A2 _3488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_58_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_58_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_73_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8215__I _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8561__A2 _3652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6572__A1 _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5127__A2 _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6875__A2 _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5678__A3 _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7824__A1 _2871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4638__A1 _4215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8001__A1 _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7964__I _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8552__A2 _3610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5620_ _0921_ as2650.stack\[5\]\[2\] _0913_ _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5366__A2 _4142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5551_ _0853_ _0854_ _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5484__I _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8304__A2 _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8270_ _3287_ _3373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5118__A2 _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5482_ _4494_ _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8855__A3 _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7221_ as2650.addr_buff\[3\] _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6866__A2 _2019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8728__C _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7152_ _2309_ _2310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7815__A1 _2774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6103_ _1375_ _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7083_ _0925_ _2256_ _2262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_140_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7204__I _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6034_ _1303_ _1306_ _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8240__A1 _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7043__A2 _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7985_ _4244_ _3107_ _3109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_54_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8791__A2 _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6936_ _2141_ _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7079__C _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6867_ _1156_ _1938_ _2077_ _0101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8543__A2 _3624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8606_ _3046_ _3697_ _3698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5818_ _1076_ _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6554__A1 _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5357__A2 _4505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6798_ _2007_ _2010_ _2011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7897__A4 _3021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8537_ as2650.addr_buff\[1\] _2538_ _3632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5749_ _1016_ _1023_ _1031_ _0029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_108_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5109__A2 _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8468_ _2825_ _0674_ _3565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_136_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7419_ _4529_ _0292_ _2556_ _2557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_8399_ _1579_ _2762_ _3498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7542__C _2340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6609__A2 _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7282__A2 _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5293__A1 _4155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5832__A3 _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8231__A1 _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7034__A2 _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8782__A2 _3525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6793__A1 _1757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5596__A2 _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6793__B2 _4520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8534__A2 _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6545__A1 _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5348__A2 _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8298__A1 _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8548__C _3331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5520__A2 _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7024__I _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5659__I0 _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6076__A3 _4174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8470__A1 _1604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9014__A3 _3216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7025__A2 _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7770_ _2386_ _2886_ _2900_ _2901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5587__A2 _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4982_ _4346_ _0292_ _4412_ _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6721_ _4195_ _1164_ _1935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_3_wb_clk_i clknet_3_2_0_wb_clk_i clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_71_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6652_ as2650.r0\[2\] _1809_ _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5603_ _0861_ _0906_ _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9371_ _0264_ clknet_leaf_76_wb_clk_i as2650.r123\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6583_ _1808_ _1813_ _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_121_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8322_ as2650.pc\[2\] _0909_ as2650.pc\[0\] _3423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__6103__I _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5534_ _4532_ _0834_ _0838_ _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8739__B _3824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8253_ _0911_ _3301_ _3356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5465_ _0770_ _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7204_ _1682_ _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8184_ _3287_ _3288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5511__A2 _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5396_ _0296_ _0662_ _0702_ _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4558__I _4138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7135_ _0924_ _2298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8461__A1 _3333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7264__A2 _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7066_ _2139_ _1905_ _2248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6017_ _0685_ _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8193__C _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5027__A1 _4420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8764__A2 _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7968_ _2160_ _3093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_42_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6919_ _2124_ _2126_ _2127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_74_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7899_ _2662_ _3023_ _3025_ _2476_ _3026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_51_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6527__A1 _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9345__CLK clknet_leaf_52_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6013__I _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6948__I _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_41_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7272__C _2411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5073__B _4408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_73_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_73_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7255__A2 _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8452__A1 _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5266__A1 _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8204__A1 _3093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7007__A2 _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8755__A2 _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5569__A2 _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8831__C _3910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8507__A2 _2539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_80_wb_clk_i_I clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7191__A1 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7019__I _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5741__A2 _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9381__D _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5250_ _0556_ _0557_ _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_114_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5181_ _0487_ _0464_ _0488_ _4502_ _0489_ _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_64_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7910__C _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9218__CLK clknet_leaf_56_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8994__A2 _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8940_ as2650.r123\[2\]\[0\] _3989_ _3990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_49_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8871_ _3939_ _3940_ _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8746__A2 _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7822_ _2948_ _2949_ _2950_ _2951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7403__C1 _2537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6757__A1 _4519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9368__CLK clknet_leaf_65_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7753_ net36 _2884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4965_ _4206_ _4543_ _4544_ _4545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_75_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6704_ _1923_ _1925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6509__A1 _4541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7684_ _2783_ _2816_ _2817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5980__A2 _4428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4896_ _4476_ _4477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6635_ _1833_ _1858_ _1864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9354_ _0247_ clknet_leaf_59_wb_clk_i as2650.stack\[7\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6566_ _1775_ _1790_ _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8305_ _2509_ _3405_ _3406_ _3407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5517_ _0799_ _0741_ _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_9285_ _0178_ clknet_leaf_27_wb_clk_i net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6497_ _1731_ _1732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5672__I _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8236_ net6 _4281_ _3339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7092__C _2243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7485__A2 _2618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5448_ _0753_ _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8682__A1 _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8167_ _3264_ _3271_ _3151_ _3272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_120_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5379_ _0354_ _4506_ _0370_ _0542_ _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_43_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8434__A1 _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7237__A2 _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7118_ _2147_ _2281_ _2283_ as2650.stack\[3\]\[0\] _2278_ _2284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_8098_ _1348_ _3209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_102_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5248__A1 _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8985__A2 _2438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7049_ as2650.r123_2\[3\]\[2\] _2237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5799__A2 _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8737__A2 _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6748__A1 as2650.r0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_8_wb_clk_i_I clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8651__C _3373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output16_I net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5420__A1 _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8223__I _2408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5971__A2 _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5723__A2 _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8673__A1 _3219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8673__B2 _3760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5487__A1 _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8425__A1 _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5239__A1 _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8976__A2 _3163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4926__I _4505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8728__A2 _1749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6739__A1 as2650.r0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7936__B1 _3061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8561__C _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4750_ _4257_ _4331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5962__A2 _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4681_ _4248_ _4261_ _4262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7164__A1 _2285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6420_ as2650.stack\[2\]\[10\] _1664_ _1667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8900__A2 _4272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6911__A1 _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6351_ _1147_ _1393_ _0505_ _0597_ _1578_ _1601_ _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_66_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5302_ _4351_ _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_143_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7467__A2 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9070_ _3770_ _3268_ _4062_ _4104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6282_ _4328_ _1360_ _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8021_ _3138_ _0549_ _3130_ _3139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_102_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5233_ _0495_ _0497_ _0501_ _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_102_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7219__A2 _2363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5164_ _4279_ _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_9_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4836__I _4170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8967__A2 _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7212__I as2650.addr_buff\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5095_ _0403_ _0307_ _0404_ _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__9190__CLK clknet_leaf_65_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8923_ _0981_ _1939_ _3976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8719__A2 _2592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8854_ _3926_ _3927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7805_ _2913_ _2934_ _2935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8785_ _3780_ _3867_ _3868_ _3869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5667__I _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5997_ _4543_ _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XPHY_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5402__B2 _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4571__I _4151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7736_ _0835_ _0827_ _2798_ _2802_ _2826_ _2867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_4948_ net7 _4528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5953__A2 _4157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7667_ _0682_ _2800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4879_ _4459_ _4460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6618_ _1845_ _1846_ _1847_ _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_53_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7598_ _0594_ _0613_ _2732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5705__A2 _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6498__I _1732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6549_ _4147_ _0540_ _1780_ _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_9337_ _0230_ clknet_leaf_77_wb_clk_i as2650.r0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8655__A1 _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9268_ _0161_ clknet_leaf_52_wb_clk_i as2650.stack\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5469__A1 _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8219_ as2650.stack\[3\]\[0\] _1918_ _1902_ as2650.stack\[0\]\[0\] as2650.stack\[1\]\[0\]
+ _1654_ _3323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
X_9199_ _0092_ clknet_leaf_47_wb_clk_i as2650.stack\[0\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8407__A1 _2694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4692__A2 _4272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8218__I _1637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7122__I _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6969__A1 _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7630__A2 _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8662__B _1496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4995__A3 _4302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5577__I as2650.addr_buff\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6197__A2 _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7697__A2 _2588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5526__B _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_3_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8646__A1 _2634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7449__A2 _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8949__A2 _3992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9071__A1 _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5920_ _0639_ _1101_ _1195_ _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5851_ _4388_ _1101_ _1130_ _1110_ _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_80_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6092__B _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6188__A2 _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7385__A1 _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4802_ _4382_ _4383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_61_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8570_ _2968_ _3644_ _3663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_34_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5782_ _4377_ _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_128_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7521_ _2635_ _2654_ _2656_ _2657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7916__B _2943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4733_ _4313_ _4314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8334__B1 _3433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7452_ _2584_ _2587_ _2588_ _2589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4664_ _4243_ _4244_ _4245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6403_ _1016_ _1644_ _1652_ _0062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5436__B _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7383_ _2520_ _2521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4595_ _4172_ _4166_ _4175_ _4176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__6111__I _4387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9122_ _0015_ clknet_leaf_42_wb_clk_i as2650.stack\[5\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6334_ _1226_ _0684_ _1583_ _1590_ _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_143_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9053_ _0821_ _1431_ _4086_ _4087_ _4088_ _4089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_6265_ _4428_ _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6112__A2 _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8004_ _3124_ _0297_ _3120_ _3125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5216_ _0328_ _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6196_ _0360_ _4541_ _4405_ _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__5871__A1 _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8038__I _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5147_ _4300_ _4522_ _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__9062__A1 _4064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7999__I0 _3115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5078_ _0386_ _0356_ _0387_ _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_42_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8906_ _3963_ _3964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4977__A3 _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8837_ _3914_ _3915_ _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7376__A1 _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6179__A2 _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7376__B2 _2513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5926__A2 _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8768_ _1558_ _1547_ _3850_ _3852_ _1513_ _3853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_90_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7826__B _2744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7719_ _2491_ _2646_ _2851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_139_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8699_ _3143_ _1383_ _3080_ _3787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_139_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8876__A1 _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7117__I _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6351__A2 _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6021__I _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8657__B _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7300__A1 _4423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7851__A2 _2522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5081__B _4345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9053__A1 _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7603__A2 _4246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8800__A1 _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7367__A1 _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7119__A1 _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8316__B1 _3390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8867__A1 _2294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8619__A1 _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7471__B _2607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6050_ _1322_ _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7842__A2 _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input7_I io_in[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5001_ _0310_ _0311_ _4325_ _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6653__I0 as2650.r123\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6952_ _2153_ _0889_ _2155_ _2157_ _2158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_66_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5903_ _0683_ _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6883_ _2090_ _2092_ _2093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_35_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8622_ _4265_ _3345_ _2353_ _3712_ _3048_ _3713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5834_ _0321_ _1094_ _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8553_ _2365_ _3646_ _3647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_5765_ _4150_ _4261_ _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_37_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7504_ _2602_ _2619_ _2639_ _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4716_ _4280_ _4297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8484_ _3415_ _3563_ _3581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8858__A1 _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5696_ _0989_ _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7435_ _1357_ _2573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8322__A3 as2650.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4647_ _4223_ _4227_ _4228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7530__A1 _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6333__A2 _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7366_ _2504_ _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4578_ _4158_ _4159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9105_ _4122_ _4133_ _4134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6317_ _1570_ _1573_ _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8086__A2 _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7297_ _1314_ _2435_ _2436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5680__I _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9036_ _4072_ _1290_ _1520_ _4073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6248_ _1492_ _1495_ _1496_ _1505_ _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_83_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4647__A2 _4227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9035__A1 _4430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6179_ _0721_ _0795_ _1436_ _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_57_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7597__A1 _2727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8794__B1 _3184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9101__B _3619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7400__I _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5072__A2 _4388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7349__A1 _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8546__B1 _3317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_27_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_27_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_71_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7275__C _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7521__A1 _2635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7824__A2 _2869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5835__A1 _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4638__A2 _4218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9026__A1 _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9251__CLK clknet_leaf_63_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8001__A2 _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9384__D _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5550_ _4488_ _4429_ _4424_ _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_30_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5481_ as2650.r123\[0\]\[7\] _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_129_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7220_ _0376_ _2358_ _2367_ _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_126_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7151_ _0857_ _2248_ _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_141_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6102_ _1374_ _4266_ _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_98_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7082_ _2183_ _2252_ _2253_ as2650.stack\[1\]\[3\] _2254_ _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_140_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5826__A1 _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6033_ _4238_ _0886_ _1304_ _1305_ _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9017__A1 _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7291__A3 _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7579__A1 _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8240__A2 _1681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7984_ _4265_ _2824_ _3108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6935_ _0967_ _2140_ _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_78_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6866_ as2650.r123_2\[2\]\[3\] _2019_ _2076_ _1980_ _2077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8605_ _3194_ _3690_ _3696_ _3697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5817_ _4513_ _1097_ _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6797_ _2004_ _2008_ _2009_ _2010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__5675__I _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6554__A2 _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8051__I _3163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8536_ _3221_ _3630_ _3631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5748_ as2650.stack\[5\]\[14\] _1021_ _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_109_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7503__A1 as2650.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8467_ _2825_ _0674_ _3564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5679_ _0966_ _0968_ _0973_ as2650.r123_2\[0\]\[0\] _0974_ _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__6306__A2 _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8700__B1 _3183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_31_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7418_ _4390_ _4352_ _2556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8398_ _3393_ _3496_ _3497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_123_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7349_ _2486_ _2487_ _2488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_46_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5817__A1 _4513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9008__A1 _4463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9019_ _1517_ _1622_ _1624_ _4056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_58_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5293__A2 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7130__I _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7990__A1 _3107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7286__B _4418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7742__A1 _2334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6545__A2 _1732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8298__A2 _4517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4929__I _4508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5808__A1 _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6076__A4 _4172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8470__A2 _4370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8564__C _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9379__D _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8136__I _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6233__A1 _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4981_ _0289_ _0291_ _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7981__A1 _2551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6720_ _1059_ _1145_ _1165_ _1934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_32_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6651_ as2650.r0\[1\] _1840_ _1880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7733__A1 net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5602_ _0865_ _0903_ _0905_ _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9147__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6582_ _4294_ _1812_ _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9370_ _0263_ clknet_leaf_76_wb_clk_i as2650.r123\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8321_ _2416_ _3422_ _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5533_ _0837_ _0598_ _4231_ _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8739__C _3088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8252_ _0909_ _3301_ _3355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5464_ _0487_ _0679_ _0743_ _0571_ _0769_ _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_133_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7203_ _2352_ _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4839__I _4143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9297__CLK clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8183_ _3055_ _3284_ _3285_ _3286_ _3287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_5395_ _0285_ _0668_ _0701_ _0295_ _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_99_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7134_ _2296_ _2286_ _2287_ as2650.stack\[3\]\[3\] _2288_ _2297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_67_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7065_ _2246_ _2247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6016_ _0670_ _1289_ _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5027__A2 _4488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7967_ _2380_ _3091_ _1481_ _3092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8490__B _4476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6918_ _2106_ _2114_ _2125_ _2126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_42_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7898_ _3020_ _3024_ _3025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6849_ _0671_ _1811_ _2060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_50_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8519_ _3391_ _3613_ _3614_ _3615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_109_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4749__I _4329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7125__I _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8452__A2 _3529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6463__A1 _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5266__A2 _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6215__A1 _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_42_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_42_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_3275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7795__I _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4777__A1 _4357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6204__I _4250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7191__A2 _2340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4701__A1 _4280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5180_ _0384_ _0482_ _0483_ _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__8575__B _2369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6454__A1 _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4608__B _4188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8870_ _2298_ _3935_ _3940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5009__A2 _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7403__B1 _2535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7821_ _2899_ _2361_ _2366_ _2950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__7403__C2 _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7752_ _2467_ _2874_ _2882_ _2598_ _2883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4964_ _4422_ _4194_ _4544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_6703_ _1923_ _1924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7683_ _2814_ _2815_ _2816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6509__A2 _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4895_ _4475_ _4476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6634_ _1833_ _1858_ _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7654__B net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5193__A1 _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9353_ _0246_ clknet_leaf_44_wb_clk_i as2650.stack\[7\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6565_ _1775_ _1790_ _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8304_ _1553_ _2538_ _3406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_121_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5516_ _0636_ _0795_ _0817_ _0820_ _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_9284_ _0177_ clknet_leaf_26_wb_clk_i net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4791__I1 as2650.r123\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6496_ _1730_ _1731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8235_ _1677_ _3335_ _2926_ _3338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5447_ _4376_ _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8682__A2 _3770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5378_ _0684_ _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8166_ _3267_ _3269_ _3270_ _3271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7117_ _2282_ _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8434__A2 _2790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8097_ _3207_ _3208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6445__A1 _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5248__A2 _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7048_ _2236_ _0123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9312__CLK clknet_leaf_18_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7829__B _2957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6748__A2 _1744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8999_ _3189_ _4038_ _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_76_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5420__A2 _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5971__A3 _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8370__A1 _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6959__I _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5863__I as2650.r123_2\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8122__A1 _3209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8673__A2 _4344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5487__A2 _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7633__B1 _2766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8976__A3 _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4998__A1 _4315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5103__I as2650.holding_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7936__A1 net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6739__A2 _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7936__B2 _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5962__A3 _4489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4680_ _4250_ _4151_ _4260_ _4261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_18_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5175__A1 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5175__B2 _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6911__A2 _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6350_ _4530_ _4387_ _4526_ _1554_ _0680_ _0758_ _1607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_122_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5706__C _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8113__A1 _3220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5301_ _4501_ _0578_ _0608_ _0285_ _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_142_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6281_ _1383_ _0754_ _0481_ _1538_ _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_115_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5232_ as2650.r123\[0\]\[4\] _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8020_ _3135_ _3137_ _3138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5163_ _0411_ _0460_ _0468_ _4225_ _0471_ _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_69_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6427__A1 _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7624__B1 _2688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9335__CLK clknet_leaf_80_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5094_ _0297_ _4331_ _0298_ _0303_ _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_69_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8922_ _3974_ _3975_ _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4989__A1 _4279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7649__B _2781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8853_ _2212_ _3899_ _3926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7927__A1 _4491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7804_ _2890_ _2902_ _2934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8324__I _3424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8784_ _1628_ _1537_ _3868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5996_ _4201_ _1268_ _1269_ _1237_ _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_80_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7735_ as2650.addr_buff\[0\] _2866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4947_ _4526_ _4527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5953__A3 _4278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7666_ _0682_ _0667_ _2799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__8352__A1 _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4878_ _4456_ _4458_ _4459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6617_ as2650.r0\[4\] _1745_ _1847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5166__A1 _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7597_ _2727_ _2730_ _2731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_88_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9336_ _0229_ clknet_3_0_0_wb_clk_i as2650.r0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6548_ _4146_ as2650.r123_2\[0\]\[4\] _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8104__A1 _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8655__A2 _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9267_ _0160_ clknet_leaf_54_wb_clk_i as2650.stack\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6479_ _1714_ _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5469__A2 _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8218_ _1637_ _3322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9198_ _0091_ clknet_leaf_46_wb_clk_i as2650.stack\[0\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8149_ _3208_ _2484_ _3249_ _3255_ _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__8407__A2 _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6418__A1 _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6969__A2 _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7091__A1 _2200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6019__I _4443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8662__C _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8591__A1 _2995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6197__A3 _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_15_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8343__A1 _3293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5157__A1 _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9208__CLK clknet_leaf_77_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9065__I _4072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8646__A2 _3727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9358__CLK clknet_leaf_59_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7082__A1 _2183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7909__A1 _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5850_ _0372_ _1103_ _1127_ _1129_ _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_73_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6092__C _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8582__A1 _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6188__A3 _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7385__A2 _4418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4801_ as2650.r0\[1\] _4382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5396__A1 _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5781_ _1062_ _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7520_ _0928_ _2655_ _2656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4732_ _4159_ _4179_ _4313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8334__A1 _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8334__B2 _2352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5148__A1 _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7451_ _4246_ _2588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4663_ as2650.idx_ctrl\[0\] _4244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8885__A2 _3949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6402_ as2650.stack\[3\]\[14\] _1642_ _1652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7382_ _2464_ _2520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4594_ _4174_ _4168_ _4175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_9121_ _0014_ clknet_leaf_39_wb_clk_i as2650.stack\[5\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6333_ as2650.psu\[3\] _1585_ _1588_ net27 _1589_ _4392_ _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XFILLER_143_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6648__A1 as2650.r0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8747__C _3765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9052_ _0732_ _0739_ _4088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6264_ _1520_ _0681_ _1521_ _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5215_ _0523_ _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8003_ _3122_ _3123_ _3124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4847__I _4197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6195_ _0394_ _1452_ _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7223__I _2357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5146_ _0448_ _0454_ _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7999__I1 _4291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5077_ _4359_ _4525_ _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7379__B _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8905_ _1390_ _3960_ _3958_ _3963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8836_ _2294_ _3912_ _3915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7376__A2 _2496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8573__A1 _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6179__A3 _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8767_ _3851_ _0593_ _1541_ _3852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7893__I as2650.addr_buff\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5979_ _1238_ _4136_ _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7718_ _2618_ _2849_ _2850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8698_ _4513_ _0292_ _3785_ _3786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_127_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5139__A1 _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7649_ _2777_ _2780_ _2781_ _2782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_60_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9319_ _0212_ clknet_3_6_0_wb_clk_i as2650.pc\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_109_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7300__A2 _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4757__I _4226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7133__I _2182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9053__A2 _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8261__B1 _3362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8800__A2 _3766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7289__B _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7367__A2 _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8564__A1 _3458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8316__A1 _3336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8316__B2 _3369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8867__A2 _3935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8619__A2 _3709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5550__A1 _4488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8567__C _3526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5000_ _4302_ _4326_ _0305_ _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5853__A2 _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__9044__A2 _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6653__I1 as2650.r123_2\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6951_ _2156_ _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_54_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5902_ _0712_ _1117_ _1178_ _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_6882_ _2058_ _2069_ _2091_ _2092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7358__A2 _2487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8555__A1 _2969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8621_ _1008_ _1544_ _3712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5833_ _0292_ _1057_ _1113_ _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_90_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8552_ _2952_ _3610_ _3646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8307__A1 _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5764_ _4223_ _1045_ _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_124_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7503_ as2650.pc\[2\] _0373_ _2639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4715_ _4295_ _4198_ _4296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8483_ _3293_ _3569_ _3579_ _3580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5695_ _0988_ _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7218__I _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7434_ _2480_ _2537_ _2567_ _1337_ _2571_ _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_120_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4646_ _4181_ _4224_ _4226_ _4227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__7662__B _2794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5541__A1 _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7365_ _2153_ _2503_ _2504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_4577_ as2650.ins_reg\[6\] _4158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9104_ _3133_ _4028_ _4133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6316_ _1411_ _1457_ _1458_ _1572_ _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_89_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7296_ _4233_ _1326_ _2434_ _2435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__7294__A1 _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9035_ _4430_ _1527_ _4072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6247_ _1499_ _1502_ _1503_ _1504_ _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_77_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9035__A2 _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8493__B _3376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6178_ _0641_ _1435_ _0722_ _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5129_ _4446_ _0436_ _0437_ _0438_ _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_84_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8794__A1 _3838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4804__B1 _4286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7349__A2 _2487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8546__A1 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8546__B2 _3624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8819_ _2208_ _3899_ _3900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_81_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_60_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_67_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_67_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7521__A2 _2654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6967__I _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7999__S _3120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7285__A1 _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6088__A2 _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7798__I _2927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7037__A1 _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8785__A1 _3780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8537__A1 as2650.addr_buff\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4950__I _4529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5267__B _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5480_ _0715_ _4440_ _0785_ _0006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7150_ _2306_ _2308_ _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6101_ _1323_ _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6079__A2 _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7081_ _2259_ _2260_ _0132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_141_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5826__A2 _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6032_ _4252_ _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_98_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7028__A1 _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7579__A2 _2553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8776__A1 _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8240__A3 _3342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7983_ _2407_ _3105_ _2434_ _3106_ _3107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__6787__B1 _1764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6934_ _2139_ _1640_ _2140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_70_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_78_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6865_ _2051_ _2075_ _2076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_126_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7200__A1 _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8604_ _3692_ _3694_ _3695_ _3696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4860__I _4406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7376__C _2514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7200__B2 _2349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5816_ _1096_ _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_91_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6796_ _0498_ _1811_ _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_22_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5357__A4 _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8535_ _1336_ _2936_ _3629_ _3630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5747_ _1012_ _1023_ _1030_ _0028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5762__A1 _4180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8466_ _3562_ _3563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5678_ as2650.r123\[0\]\[0\] _4153_ _0855_ _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_136_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7503__A2 _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8700__A1 _3219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8700__B2 _3786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7417_ _2468_ _2555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4629_ _4207_ _4209_ _4210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5691__I _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8397_ _3495_ _3496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_89_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7348_ _0863_ _4391_ _2487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_137_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7279_ _2417_ _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9018_ _4049_ _4054_ _4055_ _3742_ _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_131_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7411__I _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8767__A1 _3851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output39_I net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6027__I _4438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8519__A1 _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5866__I _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8242__I _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5753__A1 _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5505__A1 _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9006__C _3230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8455__B1 _3386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8618__S _3353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8845__C _3910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8470__A3 _3566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4945__I _4524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6769__B1 _1942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6233__A2 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7430__A1 _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4980_ _4348_ _0288_ _4506_ _0290_ _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_64_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5776__I _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5992__A1 _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6650_ _1875_ _1878_ _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_108_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8930__A1 _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5601_ as2650.stack\[5\]\[0\] _0904_ _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6581_ _1811_ _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8320_ _2178_ _3377_ _3421_ _3422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5532_ _0836_ _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_121_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8251_ _1681_ _3353_ _3354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5463_ _0384_ _0746_ _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7202_ _0877_ _1260_ _2352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8182_ _3052_ _3069_ _3071_ _3286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_5394_ _4354_ _0696_ _0699_ _0700_ _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_132_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7133_ _2182_ _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8997__A1 _4027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7064_ _2148_ _1905_ _2162_ _2246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_113_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6015_ _1288_ _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6275__C _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8749__A1 _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7421__A1 _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7966_ net51 _3090_ _3091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6917_ _2111_ _2113_ _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5983__A1 _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7897_ _2998_ _2876_ _2878_ _3021_ _3024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_23_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5686__I _4415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8062__I _4241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6848_ _0499_ _2005_ _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8921__A1 _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6779_ _1990_ _1991_ _1992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8518_ _3257_ _3596_ _3602_ _2550_ _2928_ _3614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_104_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7488__A1 _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7488__B2 _2550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8449_ _3458_ _3530_ _3544_ _3126_ _3546_ _3547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__9241__CLK clknet_leaf_55_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6160__A1 _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8988__A1 _2634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6463__A2 _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4765__I _4345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5266__A3 _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7141__I _2196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6215__A2 _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6980__I _2182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_11_wb_clk_i clknet_3_2_0_wb_clk_i clknet_leaf_11_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_122_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7479__A1 _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8428__B1 _3525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4701__A2 _4281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8979__A1 _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6454__A2 _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7403__A1 _2530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7820_ _2662_ _2871_ _2869_ _2949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7403__B2 _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9114__CLK clknet_leaf_67_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7954__A2 _3075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7751_ _2879_ _2881_ _2882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4963_ _4487_ _4543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_36_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6702_ _1922_ _1923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7682_ _2729_ _2727_ _2815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4894_ _4473_ _4474_ _4475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_71_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6633_ _1861_ _1862_ _0082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9264__CLK clknet_leaf_52_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9352_ _0245_ clknet_leaf_38_wb_clk_i as2650.stack\[7\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7654__C _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6564_ _1794_ _1795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6390__A1 _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8303_ _3401_ _3404_ _3405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5515_ _0473_ _0819_ _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_9283_ _0176_ clknet_leaf_26_wb_clk_i net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7226__I as2650.addr_buff\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6495_ as2650.r123\[0\]\[1\] as2650.r123_2\[0\]\[1\] _4145_ _1730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_69_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6130__I _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8234_ _3336_ _3335_ _3337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5446_ _0751_ _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8682__A3 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6693__A2 _1907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8165_ _0791_ _3074_ _3270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5377_ _0683_ _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8485__C _3001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7116_ _2165_ _2140_ _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8096_ _3106_ _3207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7642__A1 _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4585__I _4165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8057__I _3045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7047_ as2650.r123_2\[3\]\[1\] _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8198__A2 _3301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7829__C _2888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8998_ _2223_ _4027_ _4035_ _4037_ _4038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7949_ _1503_ _3074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_70_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5708__A1 as2650.stack\[6\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8370__A2 _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8122__A2 _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7633__A1 _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7633__B2 _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__9137__CLK clknet_leaf_46_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7936__A2 _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9287__CLK clknet_leaf_27_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8361__A2 _3428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6372__A1 _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8649__B1 _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8113__A2 _3222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5300_ _0580_ _4363_ _4501_ _0607_ _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6280_ _0744_ _1537_ _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7872__A1 _2995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5231_ _0441_ _4499_ _0539_ _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_9_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4686__A1 as2650.addr_buff\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5883__B1 _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5162_ _0461_ _4422_ _4336_ _0470_ _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_64_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7624__A1 _2757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6427__A2 _1661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7624__B2 _2736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5093_ _0303_ _0304_ _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_116_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8921_ _0616_ _3969_ _3975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8852_ _3924_ _3925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_25_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7927__A2 _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7803_ _2514_ _2932_ _2933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5938__A1 _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8783_ _3862_ _3866_ _3790_ _3867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5995_ _1236_ _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7734_ _2774_ _2864_ _2865_ _0180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4946_ _4525_ _4526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7665_ _1587_ _0748_ _2798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5964__I _4197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4877_ _4457_ _4458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6616_ as2650.r0\[5\] _1730_ _1846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5166__A2 _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6363__A1 _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7596_ _2728_ _2729_ _2730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9335_ _0228_ clknet_leaf_80_wb_clk_i as2650.r0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6547_ _1776_ _1777_ _1778_ _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__8104__A2 _4175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9266_ _0159_ clknet_leaf_54_wb_clk_i as2650.stack\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6478_ _1601_ _1051_ _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_134_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7863__A1 _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8217_ as2650.stack\[4\]\[0\] _3319_ _3320_ as2650.stack\[5\]\[0\] _4475_ _3321_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_134_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5429_ _0651_ _0732_ _0734_ _0553_ _0562_ _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_79_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9197_ _0090_ clknet_leaf_47_wb_clk_i as2650.stack\[1\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4677__A1 as2650.ins_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8148_ _3226_ _3251_ _3253_ _3254_ _3207_ _3255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_102_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8079_ _1498_ _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output21_I net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8591__A2 _3621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6197__A4 _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8250__I _3155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6106__A1 _4441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6657__A2 _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9056__B1 _3115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7606__A1 _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6409__A2 _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9030__B _2631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6373__C _1629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7909__A2 _3028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8582__A2 _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4800_ _4297_ _4380_ _4381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6188__A4 _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6593__A1 _1795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5396__A2 _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5780_ _1048_ _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7485__B _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4731_ _4183_ _4312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8334__A2 _3424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8160__I _4420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7450_ _2585_ _2586_ _2587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4662_ as2650.idx_ctrl\[1\] _4243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5148__A2 _4142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6345__A1 _1597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7542__B1 _2650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_11_wb_clk_i_I clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6401_ _1012_ _1644_ _1651_ _0061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_70_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7381_ _2416_ _2519_ _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4593_ _4173_ _4174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_116_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9120_ _0013_ clknet_leaf_38_wb_clk_i as2650.stack\[5\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6332_ _4467_ _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__9302__CLK clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6648__A2 _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9051_ _0653_ _0661_ _0732_ _0739_ _4087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_89_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6263_ _1064_ _0745_ _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4659__A1 _4238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8002_ _4542_ _1294_ _3123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5214_ _4412_ _0476_ _0522_ _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_83_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9047__B1 _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6194_ _1322_ _0447_ _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5145_ _0445_ _0453_ _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_69_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8763__C _3810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5076_ _4357_ as2650.addr_buff\[5\] _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5959__I _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8904_ _3961_ _3962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_65_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8835_ _2258_ _3908_ _3909_ as2650.stack\[6\]\[2\] _3910_ _3914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA_clkbuf_leaf_50_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8573__A2 _3648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6584__A1 _4383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8766_ _1628_ _3851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_129_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5978_ _1251_ _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7717_ _2842_ _2848_ _2849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_139_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4929_ _4508_ _4509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8697_ _2337_ _3785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7648_ _2778_ _2531_ _2534_ _1526_ _2501_ _2781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5139__A2 _4314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6336__A1 _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7579_ _0597_ _2553_ _2554_ _2713_ _2714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_125_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9318_ _0211_ clknet_leaf_30_wb_clk_i as2650.pc\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7842__C _2854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9249_ _0142_ clknet_3_1_0_wb_clk_i as2650.r123\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7064__A2 _1905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8261__B2 as2650.stack\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5075__A1 _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4773__I _4269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4822__A1 _4378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8013__A1 _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6575__A1 _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8316__A2 _3382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9325__CLK clknet_leaf_30_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4948__I net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_26_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8252__A1 _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5779__I _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6950_ _0868_ _1682_ _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_19_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5901_ _0709_ _1119_ _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_35_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6881_ _2066_ _2068_ _2091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8555__A2 _3648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8620_ _2996_ _3705_ _3711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5832_ _1060_ _1098_ _1112_ _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_62_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5613__I0 _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8551_ _2969_ _3644_ _3645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5763_ _1043_ _1044_ _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__8104__B _3214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8307__A2 _2620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7502_ _2636_ _2637_ _2638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4714_ _4294_ _4295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_8482_ _3395_ _3571_ _3563_ _3572_ _3578_ _3579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5694_ as2650.pc\[10\] _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7433_ _2486_ _2569_ _2570_ _2571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4645_ _4192_ _4225_ _4226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7364_ _0882_ _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5541__A2 _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4576_ _4156_ _4157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_9103_ as2650.psu\[3\] _4131_ _4132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6315_ _1571_ _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7234__I _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7295_ _1312_ _2433_ _2434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9034_ _1291_ _4056_ _4070_ _4071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6246_ _0867_ _4550_ _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6177_ _0567_ _0561_ _1434_ _0556_ _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_131_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8243__A1 _4531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5128_ _4493_ _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8065__I _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8794__A2 _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5059_ _0365_ _0368_ _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4804__A1 _4383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4804__B2 _4384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8546__A2 _3369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8818_ _0957_ _0427_ _3899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9348__CLK clknet_leaf_41_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8014__B _3132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8749_ _0512_ _2753_ _3757_ _3834_ _3835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_139_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6313__I _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6309__A1 _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8482__A1 _3395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7285__A2 _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8482__B2 _3572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_36_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_36_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_121_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9026__A3 _4062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8234__A1 _3336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5599__I _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8785__A2 _3867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6796__A1 _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8537__A2 _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6012__A3 _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5771__A2 _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6720__A1 _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6379__B _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6100_ _1372_ _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8473__A1 _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7080_ _0918_ _2256_ _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7989__I _2577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6031_ _4166_ _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7028__A2 _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5039__A1 _4518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8776__A2 _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7982_ _1486_ _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_66_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6787__B2 _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7938__B _3056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6933_ _0850_ _2139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6864_ _2073_ _2074_ _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_62_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7200__A2 _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8603_ _3256_ _3685_ _3691_ _2523_ _2855_ _3695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5815_ _1095_ _4268_ _1040_ _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_126_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6795_ _0362_ _1841_ _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5211__A1 _4269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6133__I _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8534_ _0979_ _1708_ _3629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5746_ as2650.stack\[5\]\[13\] _1021_ _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5762__A2 _4249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8465_ _0953_ _3561_ _3562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4789__S _4148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5677_ _0972_ _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__8700__A2 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7416_ _1308_ _2554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4628_ _4173_ _4208_ _4209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8396_ _2195_ _3494_ _3495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6711__A1 _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5514__A2 _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7347_ _2485_ _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4559_ _4139_ _4135_ _4140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_104_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8464__A1 _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7278_ net28 _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5921__B _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9017_ _1589_ _4049_ _4055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6475__B1 _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6229_ _4551_ _1271_ _0397_ _0339_ _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_131_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8767__A2 _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6308__I _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9170__CLK clknet_leaf_60_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8523__I _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6043__I _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6950__A1 _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5753__A2 _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5505__A2 _4376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5269__A1 _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7602__I _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8207__A1 _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9022__C _4058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8758__A2 _3488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6769__A1 _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7430__A2 _4390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5441__A1 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4961__I _4383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7477__C _2570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7194__A1 _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8930__A2 _3958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5600_ _0902_ _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6580_ _1810_ _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5744__A2 _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8589__B _3526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5531_ _0835_ _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_125_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8250_ _3155_ _3353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5725__C _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5462_ _0752_ _4547_ _0766_ _0767_ _0768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7201_ _2345_ _2350_ _2351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8181_ _3157_ _3163_ _1349_ _3065_ _3285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_114_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5393_ _0284_ _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7132_ _2293_ _2295_ _0148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8446__A1 _3164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7063_ _2244_ _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9193__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6014_ _1086_ _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8749__A2 _2753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6128__I _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5032__I _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7421__A2 _2553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7965_ _3089_ _3090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5432__A1 _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6916_ _0789_ _2109_ _2085_ _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_74_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7896_ _3020_ _3022_ _3023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5983__A2 _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6847_ _0788_ _2027_ _2058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8921__A2 _3969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6778_ _1961_ _1963_ _1991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8517_ _3597_ _3600_ _3596_ _3572_ _1443_ _3612_ _3613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__4943__B1 _4521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5729_ _0866_ _4466_ _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8685__A1 _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8448_ _3459_ _3545_ _3546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8379_ _3459_ _3462_ _3465_ _3478_ _3479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_105_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5207__I _4220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8437__A1 _4357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8988__A2 _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7422__I _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6215__A3 _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6482__B _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5423__A1 _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4781__I _4213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7176__A1 _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7479__A2 _2611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_51_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_51_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_127_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5117__I _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8428__A1 _3336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8428__B2 _3369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8979__A2 _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_25_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5662__A1 _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8591__C _3592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7403__A2 _2532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8600__A1 _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7750_ _2334_ _2880_ _2881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4962_ _4541_ _4542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6701_ _0866_ _1921_ _0960_ _1922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_7681_ _2786_ _2787_ _2814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4893_ _4448_ _4449_ _4474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_36_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6632_ _1201_ _1717_ _1862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5273__S0 _4196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6563_ _1725_ _1718_ _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4925__B1 _4381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9351_ _0244_ clknet_leaf_38_wb_clk_i as2650.stack\[7\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_34_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7507__I net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5193__A3 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6390__A2 _1643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8302_ _3339_ _3402_ _3403_ _3404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6411__I _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5514_ _0813_ _0565_ _0818_ _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_9282_ _0175_ clknet_leaf_26_wb_clk_i net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8667__A1 _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6494_ _1718_ _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4791__I3 as2650.r123_2\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8233_ _2387_ _3336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5445_ _0750_ _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8164_ as2650.psu\[7\] _2377_ _3268_ _3269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5376_ _0682_ _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7115_ _2280_ _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__9092__A1 _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8095_ _3190_ _3206_ _3189_ _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7242__I _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7046_ _2235_ _0122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7642__A2 _2655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8782__B _3865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5405__A1 _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8997_ _4027_ _4036_ _4037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7948_ _4490_ _2444_ _2446_ _3073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XTAP_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7879_ _2982_ _2644_ _3007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_106_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5708__A2 _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6381__A2 _4463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8658__A1 _4160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4931__A3 _4507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7861__B _2988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5892__A1 _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7152__I _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7633__A2 _2655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8692__B _3779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5644__A1 _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7149__A1 _2307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8346__B1 _1638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8897__A1 _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6372__A2 _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7327__I _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6231__I _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8649__A1 _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8649__B2 _3727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6124__A2 _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7321__A1 _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5230_ _4500_ _0524_ _0537_ _0538_ _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__7872__A2 _2996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5883__A1 _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5161_ _0469_ _0464_ _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7062__I _2243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7624__A2 _2504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5092_ _0401_ _0399_ _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_64_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5635__A1 _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8920_ _3962_ _1792_ _3964_ as2650.r123\[1\]\[4\] _3974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_42_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8851_ _3923_ _3924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_40_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7802_ _0979_ _2496_ _2931_ _2932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6406__I _1654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5399__B1 _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5994_ _1267_ _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5310__I _4426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8782_ _0341_ _3525_ _3865_ _3866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_64_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6060__A1 _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7733_ net54 _2771_ _2772_ _2865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4945_ _4524_ _4525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_36_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8888__A1 as2650.stack\[7\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7664_ _0948_ _2686_ _2796_ _2797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4876_ as2650.psu\[1\] _4457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__9381__CLK clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6615_ as2650.r0\[3\] _1762_ _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7595_ _2695_ _2717_ _2729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7560__A1 _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6363__A2 _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6546_ _1759_ _1749_ _1778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9334_ _0227_ clknet_leaf_80_wb_clk_i as2650.r0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_10_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6115__A2 _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6477_ _1084_ _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_9265_ _0158_ clknet_leaf_54_wb_clk_i as2650.stack\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7312__A1 _4220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8496__C _3592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5428_ _0654_ _0680_ _0733_ _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8216_ _1654_ _3320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7863__A2 _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9196_ _0089_ clknet_leaf_47_wb_clk_i as2650.stack\[1\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5874__A1 _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8147_ _3175_ _3226_ _3254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5359_ _0611_ _0665_ _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8078_ _3151_ _1678_ _3190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8812__A1 _3890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7029_ _2222_ _2225_ _0115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_28_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7379__A1 _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output14_I net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8879__A1 _2307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8343__A3 _3443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6051__I _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6986__I _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7303__A1 _4200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6657__A3 _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9056__A1 _1627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7606__A2 _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6409__A3 _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8803__A1 _3837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9254__CLK clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6290__A1 _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9030__C _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8567__B1 _3426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7790__A1 net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6593__A2 _1823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4730_ _4303_ _4310_ _4311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4661_ _4235_ _4241_ _4242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__7542__A1 _2661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7542__B2 _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6400_ as2650.stack\[3\]\[13\] _1642_ _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7380_ _2418_ _2466_ _2516_ _2518_ _2519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_122_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4592_ as2650.cycle\[1\] _4173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_70_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6331_ _1587_ _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_127_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9050_ _0561_ _0569_ _0653_ _0661_ _4085_ _4086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_6262_ _1519_ _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5213_ _4345_ _0485_ _0521_ _4262_ _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_8001_ _2536_ _1289_ _3122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__9047__A1 _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6193_ _1450_ _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5144_ _0449_ _0405_ _0452_ _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_96_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5075_ _0384_ _0350_ _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_96_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6281__A1 _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8903_ _3960_ _3961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8834_ _3911_ _3913_ _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6033__A1 _4238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8765_ _3843_ _3848_ _3849_ _3767_ _3850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6584__A2 _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5977_ _1250_ _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5975__I _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7716_ _2843_ _2847_ _2848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4595__A1 _4172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4928_ _4282_ _4288_ _4381_ _4385_ _4508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_142_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8696_ _3703_ _3784_ _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_90_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7647_ _2778_ _2779_ _2780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7533__A1 _2469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4859_ _4439_ _4440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6336__A2 _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9127__CLK clknet_leaf_58_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7578_ _2555_ _2712_ _2713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9317_ _0210_ clknet_leaf_25_wb_clk_i as2650.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5924__B _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6529_ _1761_ _1762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7836__A2 _2963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9248_ _0141_ clknet_leaf_63_wb_clk_i as2650.r123\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9038__A1 _3851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5215__I _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9179_ _0072_ clknet_leaf_9_wb_clk_i as2650.ins_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8526__I _3288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7064__A3 _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8261__A2 _3361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5075__A2 _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6046__I _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4822__A2 _4388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8013__A2 _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7586__B _2570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5885__I _4228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4586__A1 _4163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7524__A1 _2638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8721__B1 _3183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5838__A1 _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9029__A1 _4365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8252__A2 _3301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6263__A1 _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5900_ as2650.r123_2\[0\]\[5\] _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6880_ _2079_ _2089_ _2090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5831_ _4542_ _1099_ _1111_ _1059_ _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_61_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7763__A1 _2729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8960__B1 _3989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8550_ as2650.pc\[9\] as2650.pc\[8\] _3594_ _3644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_5762_ _4180_ _4249_ _4341_ _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_50_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7501_ _0926_ _1584_ _2637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_37_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4713_ _4285_ _4294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_6_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_6_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_124_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8481_ _2645_ _3574_ _3577_ _3076_ _3578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__7515__A1 _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5693_ _0963_ _0985_ _0987_ _0017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_33_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7432_ _1344_ _2570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4644_ _4159_ _4179_ _4225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7363_ _2501_ _2502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4575_ _4155_ _4156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9102_ _3132_ _4121_ _4131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6314_ _1532_ _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7294_ _1355_ _2432_ _2433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6245_ _4442_ _1241_ _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_9033_ _1476_ _4064_ _4065_ _4069_ _4070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_115_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8618__I1 _3705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6176_ _0442_ _0467_ _1433_ _0445_ _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_83_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5127_ _0361_ _0342_ _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8243__A2 _3345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6254__A1 _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5058_ _4297_ _0366_ _0367_ _4521_ _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_38_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4804__A2 _4140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6006__A1 _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8817_ _3837_ _3897_ _3898_ _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_38_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4823__B _4403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8748_ _1556_ _3780_ _2629_ _3833_ _3834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_71_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7506__A1 _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8679_ _0618_ _3326_ _3768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6309__A2 _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4740__A1 _4320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7285__A3 _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5296__A2 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8219__C1 as2650.stack\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4784__I _4320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8234__A2 _3335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_76_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_76_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_62_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6245__A1 _4442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8785__A3 _3868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6796__A2 _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7993__A1 _3113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6548__A2 as2650.r123_2\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4559__A1 _4139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8170__A1 _3236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9036__B _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6720__A2 _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5056__S _4516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6030_ as2650.cycle\[7\] _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input5_I io_in[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4694__I _4274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5039__A2 _4523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6236__A1 _4544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7981_ _2551_ _3104_ _3105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7984__A1 _4265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6787__A2 _1749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6932_ _4295_ _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_39_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_78_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6863_ _2052_ _2053_ _2072_ _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8602_ _3082_ _3686_ _3693_ _1276_ _3676_ _3694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_23_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5814_ _4233_ _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7200__A3 _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6794_ _1880_ _2004_ _2006_ _1969_ _2007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_50_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8533_ _3620_ _3597_ _3628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_50_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5745_ _1006_ _1023_ _1029_ _0027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5762__A3 _4341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8464_ _0945_ _2194_ _3494_ _3561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_5676_ _0294_ _0969_ _0971_ _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__8161__A1 _3265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7415_ _2469_ _2553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4627_ as2650.cycle\[0\] _4208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8395_ _0933_ _0927_ _3423_ _3494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__7245__I _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5514__A3 _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7346_ _2484_ _1311_ _2485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4558_ _4138_ _4139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_104_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8464__A2 _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7277_ _2415_ _2416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_103_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6475__A1 _4328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9016_ _3492_ _4051_ _4052_ _4053_ _4054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6475__B2 _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6228_ _1034_ _1486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_131_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8076__I _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6159_ as2650.stack\[4\]\[10\] _1420_ _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_58_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6227__A1 _1476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9315__CLK clknet_leaf_24_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7975__A1 _3088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7975__B2 _2923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7727__A1 _2854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6950__A2 _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8152__A1 _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7155__I _2312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6994__I _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput40 net40 io_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__8455__A2 _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6466__A1 _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5831__C _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8207__A2 _3310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6218__A1 _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7966__A1 net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6769__A2 _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7758__C _2888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7718__A1 _2618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8915__B1 _3967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7194__A2 _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8391__A1 _3210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5530_ net3 _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_121_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5461_ _0517_ _0593_ _4546_ _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7065__I _2246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8694__A2 _3763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7200_ _2156_ _1310_ _2346_ _2347_ _2349_ _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_133_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8180_ _3073_ _3278_ _3283_ _3284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5392_ _0486_ _0698_ _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7131_ _2294_ _2291_ _2295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6457__A1 _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7062_ _2243_ _2244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__9338__CLK clknet_leaf_39_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6013_ _1229_ _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5313__I _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6209__A1 _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7964_ _1275_ _3089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5432__A2 _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6915_ _2107_ _2114_ _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_70_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7709__A1 _2720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7895_ _2998_ _2871_ _2868_ _3021_ _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_63_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6846_ _2055_ _2056_ _2057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8382__A1 as2650.stack\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6777_ _1953_ _1962_ _1990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8516_ _3598_ _3606_ _3611_ _3070_ _3612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_17_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4943__A1 _4520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5728_ _0977_ _1016_ _1017_ _0022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4943__B2 _4522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8447_ _0946_ _3511_ _3545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_100_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8685__A2 _3773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5659_ _0951_ _0955_ _0860_ _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_87_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6696__A1 _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8378_ _3472_ _3477_ _3478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8437__A2 _3345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7329_ _4349_ _4347_ _2468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6319__I _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7948__A1 _4490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6482__C _4202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6620__A1 _4520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5423__A2 _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8373__A1 _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6989__I _2190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4934__A1 _4305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8125__A1 _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8202__C _4161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6439__A1 _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_20_wb_clk_i clknet_3_3_0_wb_clk_i clknet_leaf_20_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_111_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5111__A1 _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5662__A2 _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8061__B1 _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7488__C _2624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_30_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4961_ _4383_ _4541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6700_ _1920_ _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7680_ _2805_ _2812_ _1311_ _2813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_44_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8364__A1 _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4892_ _4448_ _4450_ _4473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6631_ as2650.r123_2\[1\]\[6\] _1729_ _1860_ _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5273__S1 _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9350_ _0243_ clknet_leaf_36_wb_clk_i as2650.stack\[7\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6562_ _1174_ _1715_ _1793_ _0080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4925__B2 _4385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8116__A1 _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8112__C _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8301_ _2581_ _4380_ _3403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5513_ _0799_ _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_9281_ _0174_ clknet_leaf_26_wb_clk_i net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8667__A2 _1476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6493_ _1713_ _1715_ _1728_ _0076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6678__A1 _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8232_ _3334_ _3335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5444_ _0672_ _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__9160__CLK clknet_leaf_58_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5350__A1 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8163_ _4176_ _1510_ _3268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5375_ net1 _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5350__B2 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7114_ _2148_ _1640_ _2212_ _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_99_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8094_ _3201_ _3205_ _4201_ _3206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_59_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9092__A2 _4028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7045_ as2650.r123_2\[3\]\[0\] _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6850__A1 _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5978__I _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8996_ _3230_ _4029_ _4036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7947_ _3069_ _3071_ _3072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7878_ _2990_ _3005_ _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_54_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5169__A1 _4304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6829_ _2037_ _2040_ _2041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_51_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8107__A1 _3211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8107__B2 _3216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8658__A2 _3265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5218__I _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4931__A4 _4510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7861__C _2888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8529__I _3623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5341__A1 _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6049__I _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8692__C _3780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7149__A2 _2291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8346__A1 as2650.stack\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8897__A2 _3949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6512__I _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9183__CLK clknet_leaf_74_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8649__A2 _3327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7321__A2 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4967__I _4546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7343__I _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5883__A2 _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5160_ _4191_ _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_123_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7085__A1 _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5091_ as2650.holding_reg\[2\] _0400_ _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5635__A2 _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8850_ _0857_ _2314_ _3923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_65_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7388__A2 _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8585__A1 _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7801_ _2926_ _2928_ _2929_ _2930_ _2931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__8585__B2 _2524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8781_ _3769_ _1812_ _3864_ _3847_ _1623_ _3865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_92_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5993_ _4174_ _4167_ _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_52_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6060__A2 _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7732_ _2205_ _2580_ _2863_ _2864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4944_ _4518_ _4523_ _4524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_80_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7663_ _2632_ _2795_ _2796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4875_ as2650.psu\[0\] _4456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_71_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6422__I _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6614_ _1839_ _1842_ _1843_ _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7594_ _2188_ _0596_ _2728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7560__A2 _2694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9333_ _0226_ clknet_leaf_80_wb_clk_i as2650.r0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6545_ _0363_ _1732_ _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5038__I _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9264_ _0157_ clknet_leaf_52_wb_clk_i as2650.stack\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6476_ _1712_ _0075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7312__A2 _2406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8215_ _1902_ _3319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5323__A1 _4477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5427_ _0730_ _0548_ _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6520__B1 _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9195_ _0088_ clknet_leaf_47_wb_clk_i as2650.stack\[1\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7253__I _4176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8146_ _2484_ _3252_ _3253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_99_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5358_ _0589_ _0664_ _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_138_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8793__B _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7076__A1 _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8077_ _3152_ _3188_ _3189_ _0199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8812__A2 _3893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5289_ _0596_ _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_75_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6823__A1 _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7028_ _0908_ _2224_ _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_60_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7379__A2 _2517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8576__A1 _2998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8979_ _1278_ _1242_ _1716_ _4018_ _4019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_128_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6339__B1 _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8879__A2 _3935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7303__A2 _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7163__I _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9056__A2 _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8264__B1 _3322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8803__A2 _3884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8208__B _3058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6290__A2 _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5411__I _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8567__A1 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8567__B2 _3652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8319__A1 _3379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7790__A2 _2885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7338__I _2476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6242__I _4208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4660_ _4237_ _4240_ _4241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__7542__A2 _2677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4591_ _4163_ _4172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6330_ _1586_ _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_122_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5305__A1 _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6502__B1 _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6261_ _1043_ _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5305__B2 _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7073__I _2243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8000_ _3121_ _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4659__A3 _4165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5212_ _0486_ _0491_ _0520_ _4247_ _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_142_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6192_ _1374_ _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__9047__A2 _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5143_ _0398_ _0451_ _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6805__A1 _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5074_ _4503_ _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8902_ _4153_ _4491_ _3960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6281__A2 _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8558__A1 _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8833_ _2290_ _3912_ _3913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_71_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7230__A1 _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8764_ _1520_ _0372_ _3849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5976_ _4417_ _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7715_ _2783_ _2789_ _2847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5792__A1 _4392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4927_ _4506_ _4507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8695_ _4441_ _3758_ _3783_ _3784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6152__I _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7646_ _2757_ _2747_ _2779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4858_ _4416_ _4437_ _4273_ _4438_ _4439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__7533__A2 _2668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6336__A3 _1592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7577_ _1580_ _0614_ _2711_ _2712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_4789_ as2650.r123\[2\]\[7\] as2650.r123_2\[2\]\[7\] _4148_ _4370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9316_ _0209_ clknet_3_2_0_wb_clk_i as2650.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6528_ as2650.r123\[0\]\[3\] as2650.r123_2\[0\]\[3\] _4144_ _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_88_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7297__A1 _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9247_ _0140_ clknet_leaf_62_wb_clk_i as2650.r123\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8079__I _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6459_ _1554_ _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9178_ _0071_ clknet_leaf_73_wb_clk_i as2650.ins_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_47_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8129_ _0687_ _2658_ _3178_ _3238_ _3239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_102_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6528__S _4144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8797__A1 _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6327__I net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6024__A2 _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5783__A1 _4220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7158__I _2315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6062__I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8021__I0 _3138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8721__A1 _3219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8721__B2 _3806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5535__A1 _4320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7288__A1 _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9221__CLK clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5838__A2 _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9029__A2 _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5850__B _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8717__I _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7621__I _2754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9371__CLK clknet_leaf_76_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9041__C _3742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6263__A2 _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5471__B1 _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5830_ _1100_ _1101_ _1109_ _1110_ _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5223__B1 _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7763__A2 _2727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8960__A1 _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5761_ _0876_ _0688_ _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7068__I _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7500_ _2181_ _0506_ _2636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_128_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4712_ _4292_ _4293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_72_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8480_ _2526_ _3562_ _3576_ _1509_ _2481_ _3577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5692_ as2650.stack\[6\]\[9\] _0986_ _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7515__A2 _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8712__A1 _3199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7431_ _2568_ _2544_ _2569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_30_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5526__A1 _4408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4643_ _4156_ _4224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_129_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6700__I _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7362_ _2396_ _1684_ _2501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4574_ as2650.ins_reg\[4\] _4155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9101_ _4128_ _4130_ _3619_ _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6313_ _1569_ _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7293_ _4169_ _4237_ _2432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5316__I _4460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9032_ _1163_ _4066_ _4068_ _4069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6244_ _1500_ _1501_ _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6175_ _0449_ _1432_ _0452_ _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8779__A1 as2650.psl\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5126_ _0432_ _0435_ _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6254__A2 _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5057_ as2650.r123\[1\]\[3\] as2650.r123\[0\]\[3\] as2650.r123_2\[1\]\[3\] as2650.r123_2\[0\]\[3\]
+ _4139_ _4516_ _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__5051__I _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5462__B1 _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5986__I _4393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6006__A2 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8816_ _1411_ _3856_ _1634_ _3898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_26_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8747_ _3790_ _0694_ _3832_ _3765_ _3833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5959_ _1232_ _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_16_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8678_ _1535_ _3767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7506__A2 _2641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7629_ _1680_ _2762_ _2763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5517__A1 _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9244__CLK clknet_leaf_39_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7706__I net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4740__A2 as2650.carry vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5226__I _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8965__C _4007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7690__A1 _2778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6493__A2 _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8219__B1 _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8219__C2 _1654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6245__A2 _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7993__A2 _3114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_45_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_72_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7745__A2 _2809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8942__A1 _4414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4559__A2 _4135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5756__A1 _4189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8221__B _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8170__A2 _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6181__A1 as2650.psl\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6720__A3 _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8473__A3 _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7433__A1 _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6236__A2 _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7980_ _3103_ _2338_ _1312_ _3104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_54_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9117__CLK clknet_leaf_41_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7984__A2 _2824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6931_ _1795_ _2136_ _2137_ _0105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_48_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6862_ _2052_ _2053_ _2072_ _2073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_35_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7736__A2 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8601_ _2372_ _2776_ _3470_ _3693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5813_ _1033_ _4261_ _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_90_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5747__A1 _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6793_ _1757_ _2005_ _1970_ _4520_ _2006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9267__CLK clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8532_ _2362_ _3626_ _3627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_91_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5744_ as2650.stack\[5\]\[12\] _1025_ _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8463_ _3559_ _3560_ _0214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8131__B _4201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5675_ _0970_ _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7526__I _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8161__A2 _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7414_ _0911_ _2528_ _2548_ _2550_ _2551_ _2552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_124_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4626_ _4163_ _4165_ _4207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5474__C _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6172__A1 _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8394_ _0933_ _3374_ _3491_ _3493_ _2415_ _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_50_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7345_ _0885_ _2484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4557_ as2650.ins_reg\[0\] _4138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7276_ _1301_ _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4885__I _4465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9015_ _3136_ _3216_ _1589_ _4053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8357__I _3456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7672__A1 _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6227_ _1476_ _1478_ _1484_ _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6475__A2 _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6158_ _0985_ _1417_ _1421_ _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_58_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7424__A1 _4529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5109_ _0397_ _0398_ _0399_ _0313_ _0417_ _0418_ _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
XTAP_3416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6089_ _4394_ _1361_ _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7727__A2 _2856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8924__A1 _3976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8820__I _3900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8152__A2 _2477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5910__A1 _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput30 net30 io_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_134_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput41 net41 io_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_107_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7663__A1 _2632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4795__I _4375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6466__A2 _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6218__A2 _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_20_wb_clk_i_I clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5620__S _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7966__A2 _3090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7718__A2 _2849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8915__A1 _3966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5729__A1 _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7194__A3 _2342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8391__A2 _3457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_117_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5460_ _4515_ _0754_ _0765_ _4538_ _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_121_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5901__A1 _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5391_ _0697_ _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_126_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7130_ _0917_ _2294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7654__A1 _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6457__A2 _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7061_ _0967_ _2166_ _2243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_113_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6012_ _1246_ _1259_ _1266_ _1285_ _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_132_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
.ends

