magic
tech gf180mcuD
magscale 1 10
timestamp 1701964108
<< metal1 >>
rect 27122 46398 27134 46450
rect 27186 46447 27198 46450
rect 27794 46447 27806 46450
rect 27186 46401 27806 46447
rect 27186 46398 27198 46401
rect 27794 46398 27806 46401
rect 27858 46447 27870 46450
rect 28354 46447 28366 46450
rect 27858 46401 28366 46447
rect 27858 46398 27870 46401
rect 28354 46398 28366 46401
rect 28418 46398 28430 46450
rect 168690 46398 168702 46450
rect 168754 46447 168766 46450
rect 169474 46447 169486 46450
rect 168754 46401 169486 46447
rect 168754 46398 168766 46401
rect 169474 46398 169486 46401
rect 169538 46398 169550 46450
rect 1344 46282 218624 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 65918 46282
rect 65970 46230 66022 46282
rect 66074 46230 66126 46282
rect 66178 46230 96638 46282
rect 96690 46230 96742 46282
rect 96794 46230 96846 46282
rect 96898 46230 127358 46282
rect 127410 46230 127462 46282
rect 127514 46230 127566 46282
rect 127618 46230 158078 46282
rect 158130 46230 158182 46282
rect 158234 46230 158286 46282
rect 158338 46230 188798 46282
rect 188850 46230 188902 46282
rect 188954 46230 189006 46282
rect 189058 46230 218624 46282
rect 1344 46196 218624 46230
rect 47742 46114 47794 46126
rect 47742 46050 47794 46062
rect 51774 46114 51826 46126
rect 51774 46050 51826 46062
rect 55806 46114 55858 46126
rect 55806 46050 55858 46062
rect 59726 46114 59778 46126
rect 59726 46050 59778 46062
rect 63534 46114 63586 46126
rect 63534 46050 63586 46062
rect 150446 46114 150498 46126
rect 150446 46050 150498 46062
rect 6974 46002 7026 46014
rect 6974 45938 7026 45950
rect 11006 46002 11058 46014
rect 11006 45938 11058 45950
rect 15038 46002 15090 46014
rect 15038 45938 15090 45950
rect 19070 46002 19122 46014
rect 19070 45938 19122 45950
rect 23102 46002 23154 46014
rect 23102 45938 23154 45950
rect 27806 46002 27858 46014
rect 27806 45938 27858 45950
rect 31614 46002 31666 46014
rect 31614 45938 31666 45950
rect 35422 46002 35474 46014
rect 35422 45938 35474 45950
rect 39230 46002 39282 46014
rect 43150 46002 43202 46014
rect 79550 46002 79602 46014
rect 40226 45950 40238 46002
rect 40290 45950 40302 46002
rect 67442 45950 67454 46002
rect 67506 45950 67518 46002
rect 71474 45950 71486 46002
rect 71538 45950 71550 46002
rect 39230 45938 39282 45950
rect 43150 45938 43202 45950
rect 79550 45938 79602 45950
rect 83582 46002 83634 46014
rect 83582 45938 83634 45950
rect 87614 46002 87666 46014
rect 87614 45938 87666 45950
rect 91646 46002 91698 46014
rect 91646 45938 91698 45950
rect 95678 46002 95730 46014
rect 95678 45938 95730 45950
rect 100158 46002 100210 46014
rect 100158 45938 100210 45950
rect 103966 46002 104018 46014
rect 103966 45938 104018 45950
rect 107774 46002 107826 46014
rect 107774 45938 107826 45950
rect 111694 46002 111746 46014
rect 111694 45938 111746 45950
rect 115502 46002 115554 46014
rect 115502 45938 115554 45950
rect 119310 46002 119362 46014
rect 119310 45938 119362 45950
rect 123902 46002 123954 46014
rect 123902 45938 123954 45950
rect 127934 46002 127986 46014
rect 127934 45938 127986 45950
rect 131966 46002 132018 46014
rect 131966 45938 132018 45950
rect 135998 46002 136050 46014
rect 135998 45938 136050 45950
rect 140030 46002 140082 46014
rect 140030 45938 140082 45950
rect 144062 46002 144114 46014
rect 144062 45938 144114 45950
rect 156158 46002 156210 46014
rect 156158 45938 156210 45950
rect 160190 46002 160242 46014
rect 160190 45938 160242 45950
rect 164222 46002 164274 46014
rect 164222 45938 164274 45950
rect 168702 46002 168754 46014
rect 168702 45938 168754 45950
rect 172510 46002 172562 46014
rect 172510 45938 172562 45950
rect 176318 46002 176370 46014
rect 176318 45938 176370 45950
rect 180238 46002 180290 46014
rect 180238 45938 180290 45950
rect 184046 46002 184098 46014
rect 184046 45938 184098 45950
rect 187854 46002 187906 46014
rect 187854 45938 187906 45950
rect 192446 46002 192498 46014
rect 196478 46002 196530 46014
rect 193106 45950 193118 46002
rect 193170 45950 193182 46002
rect 192446 45938 192498 45950
rect 196478 45938 196530 45950
rect 200510 46002 200562 46014
rect 200510 45938 200562 45950
rect 204542 46002 204594 46014
rect 208574 46002 208626 46014
rect 205202 45950 205214 46002
rect 205266 45950 205278 46002
rect 204542 45938 204594 45950
rect 208574 45938 208626 45950
rect 212606 46002 212658 46014
rect 212606 45938 212658 45950
rect 216638 46002 216690 46014
rect 217522 45950 217534 46002
rect 217586 45950 217598 46002
rect 216638 45938 216690 45950
rect 15262 45890 15314 45902
rect 7410 45838 7422 45890
rect 7474 45838 7486 45890
rect 11218 45838 11230 45890
rect 11282 45838 11294 45890
rect 15262 45826 15314 45838
rect 15822 45890 15874 45902
rect 15822 45826 15874 45838
rect 19294 45890 19346 45902
rect 19294 45826 19346 45838
rect 19854 45890 19906 45902
rect 19854 45826 19906 45838
rect 23326 45890 23378 45902
rect 23326 45826 23378 45838
rect 23886 45890 23938 45902
rect 23886 45826 23938 45838
rect 28366 45890 28418 45902
rect 28366 45826 28418 45838
rect 28926 45890 28978 45902
rect 28926 45826 28978 45838
rect 32174 45890 32226 45902
rect 32174 45826 32226 45838
rect 32734 45890 32786 45902
rect 32734 45826 32786 45838
rect 35982 45890 36034 45902
rect 35982 45826 36034 45838
rect 36542 45890 36594 45902
rect 36542 45826 36594 45838
rect 39790 45890 39842 45902
rect 39790 45826 39842 45838
rect 43598 45890 43650 45902
rect 43598 45826 43650 45838
rect 44158 45890 44210 45902
rect 55134 45890 55186 45902
rect 79774 45890 79826 45902
rect 50082 45838 50094 45890
rect 50146 45838 50158 45890
rect 54114 45838 54126 45890
rect 54178 45838 54190 45890
rect 58146 45838 58158 45890
rect 58210 45838 58222 45890
rect 62066 45838 62078 45890
rect 62130 45838 62142 45890
rect 65874 45838 65886 45890
rect 65938 45838 65950 45890
rect 69682 45838 69694 45890
rect 69746 45838 69758 45890
rect 73490 45838 73502 45890
rect 73554 45838 73566 45890
rect 44158 45826 44210 45838
rect 55134 45826 55186 45838
rect 79774 45826 79826 45838
rect 83806 45890 83858 45902
rect 83806 45826 83858 45838
rect 87838 45890 87890 45902
rect 87838 45826 87890 45838
rect 91870 45890 91922 45902
rect 91870 45826 91922 45838
rect 95902 45890 95954 45902
rect 108334 45890 108386 45902
rect 100818 45838 100830 45890
rect 100882 45838 100894 45890
rect 104626 45838 104638 45890
rect 104690 45838 104702 45890
rect 95902 45826 95954 45838
rect 108334 45826 108386 45838
rect 112142 45890 112194 45902
rect 112142 45826 112194 45838
rect 116062 45890 116114 45902
rect 116062 45826 116114 45838
rect 120094 45890 120146 45902
rect 120094 45826 120146 45838
rect 124126 45890 124178 45902
rect 124126 45826 124178 45838
rect 128158 45890 128210 45902
rect 128158 45826 128210 45838
rect 132190 45890 132242 45902
rect 156382 45890 156434 45902
rect 188638 45890 188690 45902
rect 136434 45838 136446 45890
rect 136498 45838 136510 45890
rect 140466 45838 140478 45890
rect 140530 45838 140542 45890
rect 144498 45838 144510 45890
rect 144562 45838 144574 45890
rect 152786 45838 152798 45890
rect 152850 45838 152862 45890
rect 160626 45838 160638 45890
rect 160690 45838 160702 45890
rect 164658 45838 164670 45890
rect 164722 45838 164734 45890
rect 169474 45838 169486 45890
rect 169538 45838 169550 45890
rect 173282 45838 173294 45890
rect 173346 45838 173358 45890
rect 177090 45838 177102 45890
rect 177154 45838 177166 45890
rect 180898 45838 180910 45890
rect 180962 45838 180974 45890
rect 184818 45838 184830 45890
rect 184882 45838 184894 45890
rect 132190 45826 132242 45838
rect 156382 45826 156434 45838
rect 188638 45826 188690 45838
rect 192670 45890 192722 45902
rect 192670 45826 192722 45838
rect 196702 45890 196754 45902
rect 196702 45826 196754 45838
rect 200734 45890 200786 45902
rect 200734 45826 200786 45838
rect 204766 45890 204818 45902
rect 204766 45826 204818 45838
rect 208798 45890 208850 45902
rect 212818 45838 212830 45890
rect 212882 45838 212894 45890
rect 216850 45838 216862 45890
rect 216914 45838 216926 45890
rect 208798 45826 208850 45838
rect 66558 45778 66610 45790
rect 12338 45726 12350 45778
rect 12402 45726 12414 45778
rect 66558 45714 66610 45726
rect 189198 45778 189250 45790
rect 189198 45714 189250 45726
rect 197262 45778 197314 45790
rect 197262 45714 197314 45726
rect 201294 45778 201346 45790
rect 201294 45714 201346 45726
rect 209358 45778 209410 45790
rect 213938 45726 213950 45778
rect 214002 45726 214014 45778
rect 209358 45714 209410 45726
rect 50542 45666 50594 45678
rect 7186 45614 7198 45666
rect 7250 45614 7262 45666
rect 50542 45602 50594 45614
rect 58942 45666 58994 45678
rect 58942 45602 58994 45614
rect 62750 45666 62802 45678
rect 62750 45602 62802 45614
rect 70366 45666 70418 45678
rect 70366 45602 70418 45614
rect 74174 45666 74226 45678
rect 132526 45666 132578 45678
rect 80098 45614 80110 45666
rect 80162 45614 80174 45666
rect 84130 45614 84142 45666
rect 84194 45614 84206 45666
rect 88162 45614 88174 45666
rect 88226 45614 88238 45666
rect 92194 45614 92206 45666
rect 92258 45614 92270 45666
rect 96226 45614 96238 45666
rect 96290 45614 96302 45666
rect 101042 45614 101054 45666
rect 101106 45614 101118 45666
rect 104850 45614 104862 45666
rect 104914 45614 104926 45666
rect 108658 45614 108670 45666
rect 108722 45614 108734 45666
rect 112466 45614 112478 45666
rect 112530 45614 112542 45666
rect 116386 45614 116398 45666
rect 116450 45614 116462 45666
rect 120418 45614 120430 45666
rect 120482 45614 120494 45666
rect 124450 45614 124462 45666
rect 124514 45614 124526 45666
rect 128482 45614 128494 45666
rect 128546 45614 128558 45666
rect 74174 45602 74226 45614
rect 132526 45602 132578 45614
rect 136222 45666 136274 45678
rect 136222 45602 136274 45614
rect 140254 45666 140306 45678
rect 140254 45602 140306 45614
rect 144286 45666 144338 45678
rect 144286 45602 144338 45614
rect 153246 45666 153298 45678
rect 153246 45602 153298 45614
rect 156718 45666 156770 45678
rect 156718 45602 156770 45614
rect 160414 45666 160466 45678
rect 169262 45666 169314 45678
rect 164434 45614 164446 45666
rect 164498 45614 164510 45666
rect 173058 45614 173070 45666
rect 173122 45614 173134 45666
rect 176866 45614 176878 45666
rect 176930 45614 176942 45666
rect 180674 45614 180686 45666
rect 180738 45614 180750 45666
rect 184594 45614 184606 45666
rect 184658 45614 184670 45666
rect 160414 45602 160466 45614
rect 169262 45602 169314 45614
rect 1344 45498 218624 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 50558 45498
rect 50610 45446 50662 45498
rect 50714 45446 50766 45498
rect 50818 45446 81278 45498
rect 81330 45446 81382 45498
rect 81434 45446 81486 45498
rect 81538 45446 111998 45498
rect 112050 45446 112102 45498
rect 112154 45446 112206 45498
rect 112258 45446 142718 45498
rect 142770 45446 142822 45498
rect 142874 45446 142926 45498
rect 142978 45446 173438 45498
rect 173490 45446 173542 45498
rect 173594 45446 173646 45498
rect 173698 45446 204158 45498
rect 204210 45446 204262 45498
rect 204314 45446 204366 45498
rect 204418 45446 218624 45498
rect 1344 45412 218624 45446
rect 153358 45330 153410 45342
rect 153358 45266 153410 45278
rect 140590 45218 140642 45230
rect 140590 45154 140642 45166
rect 78878 45106 78930 45118
rect 78306 45054 78318 45106
rect 78370 45054 78382 45106
rect 141586 45054 141598 45106
rect 141650 45054 141662 45106
rect 152338 45054 152350 45106
rect 152402 45054 152414 45106
rect 78878 45042 78930 45054
rect 75966 44994 76018 45006
rect 75966 44930 76018 44942
rect 135214 44994 135266 45006
rect 135214 44930 135266 44942
rect 138126 44994 138178 45006
rect 138126 44930 138178 44942
rect 138686 44994 138738 45006
rect 138686 44930 138738 44942
rect 139694 44994 139746 45006
rect 139694 44930 139746 44942
rect 139806 44994 139858 45006
rect 139806 44930 139858 44942
rect 152126 44994 152178 45006
rect 152126 44930 152178 44942
rect 1344 44714 218624 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 65918 44714
rect 65970 44662 66022 44714
rect 66074 44662 66126 44714
rect 66178 44662 96638 44714
rect 96690 44662 96742 44714
rect 96794 44662 96846 44714
rect 96898 44662 127358 44714
rect 127410 44662 127462 44714
rect 127514 44662 127566 44714
rect 127618 44662 158078 44714
rect 158130 44662 158182 44714
rect 158234 44662 158286 44714
rect 158338 44662 188798 44714
rect 188850 44662 188902 44714
rect 188954 44662 189006 44714
rect 189058 44662 218624 44714
rect 1344 44628 218624 44662
rect 132626 44382 132638 44434
rect 132690 44382 132702 44434
rect 134754 44382 134766 44434
rect 134818 44382 134830 44434
rect 135874 44382 135886 44434
rect 135938 44382 135950 44434
rect 138002 44382 138014 44434
rect 138066 44382 138078 44434
rect 139682 44382 139694 44434
rect 139746 44382 139758 44434
rect 141810 44382 141822 44434
rect 141874 44382 141886 44434
rect 131954 44270 131966 44322
rect 132018 44270 132030 44322
rect 135090 44270 135102 44322
rect 135154 44270 135166 44322
rect 138898 44270 138910 44322
rect 138962 44270 138974 44322
rect 1344 43930 218624 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 50558 43930
rect 50610 43878 50662 43930
rect 50714 43878 50766 43930
rect 50818 43878 81278 43930
rect 81330 43878 81382 43930
rect 81434 43878 81486 43930
rect 81538 43878 111998 43930
rect 112050 43878 112102 43930
rect 112154 43878 112206 43930
rect 112258 43878 142718 43930
rect 142770 43878 142822 43930
rect 142874 43878 142926 43930
rect 142978 43878 173438 43930
rect 173490 43878 173542 43930
rect 173594 43878 173646 43930
rect 173698 43878 204158 43930
rect 204210 43878 204262 43930
rect 204314 43878 204366 43930
rect 204418 43878 218624 43930
rect 1344 43844 218624 43878
rect 135886 43650 135938 43662
rect 135886 43586 135938 43598
rect 136110 43650 136162 43662
rect 139682 43598 139694 43650
rect 139746 43598 139758 43650
rect 136110 43586 136162 43598
rect 135774 43538 135826 43550
rect 135774 43474 135826 43486
rect 136222 43538 136274 43550
rect 140354 43486 140366 43538
rect 140418 43486 140430 43538
rect 136222 43474 136274 43486
rect 135102 43426 135154 43438
rect 135102 43362 135154 43374
rect 137230 43426 137282 43438
rect 137554 43374 137566 43426
rect 137618 43374 137630 43426
rect 137230 43362 137282 43374
rect 1344 43146 218624 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 65918 43146
rect 65970 43094 66022 43146
rect 66074 43094 66126 43146
rect 66178 43094 96638 43146
rect 96690 43094 96742 43146
rect 96794 43094 96846 43146
rect 96898 43094 127358 43146
rect 127410 43094 127462 43146
rect 127514 43094 127566 43146
rect 127618 43094 158078 43146
rect 158130 43094 158182 43146
rect 158234 43094 158286 43146
rect 158338 43094 188798 43146
rect 188850 43094 188902 43146
rect 188954 43094 189006 43146
rect 189058 43094 218624 43146
rect 1344 43060 218624 43094
rect 137790 42978 137842 42990
rect 137790 42914 137842 42926
rect 138126 42978 138178 42990
rect 138126 42914 138178 42926
rect 137902 42754 137954 42766
rect 137902 42690 137954 42702
rect 137790 42530 137842 42542
rect 137790 42466 137842 42478
rect 1344 42362 218624 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 50558 42362
rect 50610 42310 50662 42362
rect 50714 42310 50766 42362
rect 50818 42310 81278 42362
rect 81330 42310 81382 42362
rect 81434 42310 81486 42362
rect 81538 42310 111998 42362
rect 112050 42310 112102 42362
rect 112154 42310 112206 42362
rect 112258 42310 142718 42362
rect 142770 42310 142822 42362
rect 142874 42310 142926 42362
rect 142978 42310 173438 42362
rect 173490 42310 173542 42362
rect 173594 42310 173646 42362
rect 173698 42310 204158 42362
rect 204210 42310 204262 42362
rect 204314 42310 204366 42362
rect 204418 42310 218624 42362
rect 1344 42276 218624 42310
rect 1344 41578 218624 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 65918 41578
rect 65970 41526 66022 41578
rect 66074 41526 66126 41578
rect 66178 41526 96638 41578
rect 96690 41526 96742 41578
rect 96794 41526 96846 41578
rect 96898 41526 127358 41578
rect 127410 41526 127462 41578
rect 127514 41526 127566 41578
rect 127618 41526 158078 41578
rect 158130 41526 158182 41578
rect 158234 41526 158286 41578
rect 158338 41526 188798 41578
rect 188850 41526 188902 41578
rect 188954 41526 189006 41578
rect 189058 41526 218624 41578
rect 1344 41492 218624 41526
rect 1344 40794 218624 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 50558 40794
rect 50610 40742 50662 40794
rect 50714 40742 50766 40794
rect 50818 40742 81278 40794
rect 81330 40742 81382 40794
rect 81434 40742 81486 40794
rect 81538 40742 111998 40794
rect 112050 40742 112102 40794
rect 112154 40742 112206 40794
rect 112258 40742 142718 40794
rect 142770 40742 142822 40794
rect 142874 40742 142926 40794
rect 142978 40742 173438 40794
rect 173490 40742 173542 40794
rect 173594 40742 173646 40794
rect 173698 40742 204158 40794
rect 204210 40742 204262 40794
rect 204314 40742 204366 40794
rect 204418 40742 218624 40794
rect 1344 40708 218624 40742
rect 1344 40010 218624 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 65918 40010
rect 65970 39958 66022 40010
rect 66074 39958 66126 40010
rect 66178 39958 96638 40010
rect 96690 39958 96742 40010
rect 96794 39958 96846 40010
rect 96898 39958 127358 40010
rect 127410 39958 127462 40010
rect 127514 39958 127566 40010
rect 127618 39958 158078 40010
rect 158130 39958 158182 40010
rect 158234 39958 158286 40010
rect 158338 39958 188798 40010
rect 188850 39958 188902 40010
rect 188954 39958 189006 40010
rect 189058 39958 218624 40010
rect 1344 39924 218624 39958
rect 1344 39226 218624 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 50558 39226
rect 50610 39174 50662 39226
rect 50714 39174 50766 39226
rect 50818 39174 81278 39226
rect 81330 39174 81382 39226
rect 81434 39174 81486 39226
rect 81538 39174 111998 39226
rect 112050 39174 112102 39226
rect 112154 39174 112206 39226
rect 112258 39174 142718 39226
rect 142770 39174 142822 39226
rect 142874 39174 142926 39226
rect 142978 39174 173438 39226
rect 173490 39174 173542 39226
rect 173594 39174 173646 39226
rect 173698 39174 204158 39226
rect 204210 39174 204262 39226
rect 204314 39174 204366 39226
rect 204418 39174 218624 39226
rect 1344 39140 218624 39174
rect 1344 38442 218624 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 65918 38442
rect 65970 38390 66022 38442
rect 66074 38390 66126 38442
rect 66178 38390 96638 38442
rect 96690 38390 96742 38442
rect 96794 38390 96846 38442
rect 96898 38390 127358 38442
rect 127410 38390 127462 38442
rect 127514 38390 127566 38442
rect 127618 38390 158078 38442
rect 158130 38390 158182 38442
rect 158234 38390 158286 38442
rect 158338 38390 188798 38442
rect 188850 38390 188902 38442
rect 188954 38390 189006 38442
rect 189058 38390 218624 38442
rect 1344 38356 218624 38390
rect 1344 37658 218624 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 50558 37658
rect 50610 37606 50662 37658
rect 50714 37606 50766 37658
rect 50818 37606 81278 37658
rect 81330 37606 81382 37658
rect 81434 37606 81486 37658
rect 81538 37606 111998 37658
rect 112050 37606 112102 37658
rect 112154 37606 112206 37658
rect 112258 37606 142718 37658
rect 142770 37606 142822 37658
rect 142874 37606 142926 37658
rect 142978 37606 173438 37658
rect 173490 37606 173542 37658
rect 173594 37606 173646 37658
rect 173698 37606 204158 37658
rect 204210 37606 204262 37658
rect 204314 37606 204366 37658
rect 204418 37606 218624 37658
rect 1344 37572 218624 37606
rect 119298 37214 119310 37266
rect 119362 37214 119374 37266
rect 118750 37154 118802 37166
rect 124226 37102 124238 37154
rect 124290 37102 124302 37154
rect 118750 37090 118802 37102
rect 1344 36874 218624 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 65918 36874
rect 65970 36822 66022 36874
rect 66074 36822 66126 36874
rect 66178 36822 96638 36874
rect 96690 36822 96742 36874
rect 96794 36822 96846 36874
rect 96898 36822 127358 36874
rect 127410 36822 127462 36874
rect 127514 36822 127566 36874
rect 127618 36822 158078 36874
rect 158130 36822 158182 36874
rect 158234 36822 158286 36874
rect 158338 36822 188798 36874
rect 188850 36822 188902 36874
rect 188954 36822 189006 36874
rect 189058 36822 218624 36874
rect 1344 36788 218624 36822
rect 131058 36430 131070 36482
rect 131122 36430 131134 36482
rect 135986 36318 135998 36370
rect 136050 36318 136062 36370
rect 130510 36258 130562 36270
rect 130510 36194 130562 36206
rect 1344 36090 218624 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 50558 36090
rect 50610 36038 50662 36090
rect 50714 36038 50766 36090
rect 50818 36038 81278 36090
rect 81330 36038 81382 36090
rect 81434 36038 81486 36090
rect 81538 36038 111998 36090
rect 112050 36038 112102 36090
rect 112154 36038 112206 36090
rect 112258 36038 142718 36090
rect 142770 36038 142822 36090
rect 142874 36038 142926 36090
rect 142978 36038 173438 36090
rect 173490 36038 173542 36090
rect 173594 36038 173646 36090
rect 173698 36038 204158 36090
rect 204210 36038 204262 36090
rect 204314 36038 204366 36090
rect 204418 36038 218624 36090
rect 1344 36004 218624 36038
rect 1344 35306 218624 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 65918 35306
rect 65970 35254 66022 35306
rect 66074 35254 66126 35306
rect 66178 35254 96638 35306
rect 96690 35254 96742 35306
rect 96794 35254 96846 35306
rect 96898 35254 127358 35306
rect 127410 35254 127462 35306
rect 127514 35254 127566 35306
rect 127618 35254 158078 35306
rect 158130 35254 158182 35306
rect 158234 35254 158286 35306
rect 158338 35254 188798 35306
rect 188850 35254 188902 35306
rect 188954 35254 189006 35306
rect 189058 35254 218624 35306
rect 1344 35220 218624 35254
rect 1344 34522 218624 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 50558 34522
rect 50610 34470 50662 34522
rect 50714 34470 50766 34522
rect 50818 34470 81278 34522
rect 81330 34470 81382 34522
rect 81434 34470 81486 34522
rect 81538 34470 111998 34522
rect 112050 34470 112102 34522
rect 112154 34470 112206 34522
rect 112258 34470 142718 34522
rect 142770 34470 142822 34522
rect 142874 34470 142926 34522
rect 142978 34470 173438 34522
rect 173490 34470 173542 34522
rect 173594 34470 173646 34522
rect 173698 34470 204158 34522
rect 204210 34470 204262 34522
rect 204314 34470 204366 34522
rect 204418 34470 218624 34522
rect 1344 34436 218624 34470
rect 1344 33738 218624 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 65918 33738
rect 65970 33686 66022 33738
rect 66074 33686 66126 33738
rect 66178 33686 96638 33738
rect 96690 33686 96742 33738
rect 96794 33686 96846 33738
rect 96898 33686 127358 33738
rect 127410 33686 127462 33738
rect 127514 33686 127566 33738
rect 127618 33686 158078 33738
rect 158130 33686 158182 33738
rect 158234 33686 158286 33738
rect 158338 33686 188798 33738
rect 188850 33686 188902 33738
rect 188954 33686 189006 33738
rect 189058 33686 218624 33738
rect 1344 33652 218624 33686
rect 1344 32954 218624 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 50558 32954
rect 50610 32902 50662 32954
rect 50714 32902 50766 32954
rect 50818 32902 81278 32954
rect 81330 32902 81382 32954
rect 81434 32902 81486 32954
rect 81538 32902 111998 32954
rect 112050 32902 112102 32954
rect 112154 32902 112206 32954
rect 112258 32902 142718 32954
rect 142770 32902 142822 32954
rect 142874 32902 142926 32954
rect 142978 32902 173438 32954
rect 173490 32902 173542 32954
rect 173594 32902 173646 32954
rect 173698 32902 204158 32954
rect 204210 32902 204262 32954
rect 204314 32902 204366 32954
rect 204418 32902 218624 32954
rect 1344 32868 218624 32902
rect 117182 32786 117234 32798
rect 117182 32722 117234 32734
rect 116722 32510 116734 32562
rect 116786 32510 116798 32562
rect 112578 32398 112590 32450
rect 112642 32398 112654 32450
rect 1344 32170 218624 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 65918 32170
rect 65970 32118 66022 32170
rect 66074 32118 66126 32170
rect 66178 32118 96638 32170
rect 96690 32118 96742 32170
rect 96794 32118 96846 32170
rect 96898 32118 127358 32170
rect 127410 32118 127462 32170
rect 127514 32118 127566 32170
rect 127618 32118 158078 32170
rect 158130 32118 158182 32170
rect 158234 32118 158286 32170
rect 158338 32118 188798 32170
rect 188850 32118 188902 32170
rect 188954 32118 189006 32170
rect 189058 32118 218624 32170
rect 1344 32084 218624 32118
rect 1344 31386 218624 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 50558 31386
rect 50610 31334 50662 31386
rect 50714 31334 50766 31386
rect 50818 31334 81278 31386
rect 81330 31334 81382 31386
rect 81434 31334 81486 31386
rect 81538 31334 111998 31386
rect 112050 31334 112102 31386
rect 112154 31334 112206 31386
rect 112258 31334 142718 31386
rect 142770 31334 142822 31386
rect 142874 31334 142926 31386
rect 142978 31334 173438 31386
rect 173490 31334 173542 31386
rect 173594 31334 173646 31386
rect 173698 31334 204158 31386
rect 204210 31334 204262 31386
rect 204314 31334 204366 31386
rect 204418 31334 218624 31386
rect 1344 31300 218624 31334
rect 117294 31218 117346 31230
rect 117294 31154 117346 31166
rect 108882 30942 108894 30994
rect 108946 30942 108958 30994
rect 116722 30942 116734 30994
rect 116786 30942 116798 30994
rect 137330 30942 137342 30994
rect 137394 30942 137406 30994
rect 109454 30882 109506 30894
rect 108210 30830 108222 30882
rect 108274 30830 108286 30882
rect 109454 30818 109506 30830
rect 109902 30882 109954 30894
rect 109902 30818 109954 30830
rect 113598 30882 113650 30894
rect 136334 30882 136386 30894
rect 116050 30830 116062 30882
rect 116114 30830 116126 30882
rect 113598 30818 113650 30830
rect 136334 30818 136386 30830
rect 136782 30882 136834 30894
rect 138114 30830 138126 30882
rect 138178 30830 138190 30882
rect 140242 30830 140254 30882
rect 140306 30830 140318 30882
rect 136782 30818 136834 30830
rect 1344 30602 218624 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 65918 30602
rect 65970 30550 66022 30602
rect 66074 30550 66126 30602
rect 66178 30550 96638 30602
rect 96690 30550 96742 30602
rect 96794 30550 96846 30602
rect 96898 30550 127358 30602
rect 127410 30550 127462 30602
rect 127514 30550 127566 30602
rect 127618 30550 158078 30602
rect 158130 30550 158182 30602
rect 158234 30550 158286 30602
rect 158338 30550 188798 30602
rect 188850 30550 188902 30602
rect 188954 30550 189006 30602
rect 189058 30550 218624 30602
rect 1344 30516 218624 30550
rect 113374 30322 113426 30334
rect 135762 30270 135774 30322
rect 135826 30270 135838 30322
rect 113374 30258 113426 30270
rect 96686 30210 96738 30222
rect 104974 30210 105026 30222
rect 117630 30210 117682 30222
rect 129950 30210 130002 30222
rect 96226 30158 96238 30210
rect 96290 30158 96302 30210
rect 104402 30158 104414 30210
rect 104466 30158 104478 30210
rect 112354 30158 112366 30210
rect 112418 30158 112430 30210
rect 117954 30158 117966 30210
rect 118018 30158 118030 30210
rect 128930 30158 128942 30210
rect 128994 30158 129006 30210
rect 96686 30146 96738 30158
rect 104974 30146 105026 30158
rect 117630 30146 117682 30158
rect 129950 30146 130002 30158
rect 132638 30210 132690 30222
rect 136222 30210 136274 30222
rect 132850 30158 132862 30210
rect 132914 30158 132926 30210
rect 132638 30146 132690 30158
rect 136222 30146 136274 30158
rect 97134 30098 97186 30110
rect 105422 30098 105474 30110
rect 112926 30098 112978 30110
rect 129502 30098 129554 30110
rect 95442 30046 95454 30098
rect 95506 30046 95518 30098
rect 103730 30046 103742 30098
rect 103794 30046 103806 30098
rect 111682 30046 111694 30098
rect 111746 30046 111758 30098
rect 118738 30046 118750 30098
rect 118802 30046 118814 30098
rect 128258 30046 128270 30098
rect 128322 30046 128334 30098
rect 133634 30046 133646 30098
rect 133698 30046 133710 30098
rect 97134 30034 97186 30046
rect 105422 30034 105474 30046
rect 112926 30034 112978 30046
rect 129502 30034 129554 30046
rect 121326 29986 121378 29998
rect 121326 29922 121378 29934
rect 1344 29818 218624 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 50558 29818
rect 50610 29766 50662 29818
rect 50714 29766 50766 29818
rect 50818 29766 81278 29818
rect 81330 29766 81382 29818
rect 81434 29766 81486 29818
rect 81538 29766 111998 29818
rect 112050 29766 112102 29818
rect 112154 29766 112206 29818
rect 112258 29766 142718 29818
rect 142770 29766 142822 29818
rect 142874 29766 142926 29818
rect 142978 29766 173438 29818
rect 173490 29766 173542 29818
rect 173594 29766 173646 29818
rect 173698 29766 204158 29818
rect 204210 29766 204262 29818
rect 204314 29766 204366 29818
rect 204418 29766 218624 29818
rect 1344 29732 218624 29766
rect 101278 29650 101330 29662
rect 101278 29586 101330 29598
rect 125358 29650 125410 29662
rect 125358 29586 125410 29598
rect 133982 29650 134034 29662
rect 133982 29586 134034 29598
rect 134430 29650 134482 29662
rect 134430 29586 134482 29598
rect 135762 29486 135774 29538
rect 135826 29486 135838 29538
rect 100818 29374 100830 29426
rect 100882 29374 100894 29426
rect 124450 29374 124462 29426
rect 124514 29374 124526 29426
rect 134978 29374 134990 29426
rect 135042 29374 135054 29426
rect 101726 29314 101778 29326
rect 124910 29314 124962 29326
rect 100034 29262 100046 29314
rect 100098 29262 100110 29314
rect 123666 29262 123678 29314
rect 123730 29262 123742 29314
rect 137890 29262 137902 29314
rect 137954 29262 137966 29314
rect 101726 29250 101778 29262
rect 124910 29250 124962 29262
rect 1344 29034 218624 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 65918 29034
rect 65970 28982 66022 29034
rect 66074 28982 66126 29034
rect 66178 28982 96638 29034
rect 96690 28982 96742 29034
rect 96794 28982 96846 29034
rect 96898 28982 127358 29034
rect 127410 28982 127462 29034
rect 127514 28982 127566 29034
rect 127618 28982 158078 29034
rect 158130 28982 158182 29034
rect 158234 28982 158286 29034
rect 158338 28982 188798 29034
rect 188850 28982 188902 29034
rect 188954 28982 189006 29034
rect 189058 28982 218624 29034
rect 1344 28948 218624 28982
rect 1344 28250 218624 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 50558 28250
rect 50610 28198 50662 28250
rect 50714 28198 50766 28250
rect 50818 28198 81278 28250
rect 81330 28198 81382 28250
rect 81434 28198 81486 28250
rect 81538 28198 111998 28250
rect 112050 28198 112102 28250
rect 112154 28198 112206 28250
rect 112258 28198 142718 28250
rect 142770 28198 142822 28250
rect 142874 28198 142926 28250
rect 142978 28198 173438 28250
rect 173490 28198 173542 28250
rect 173594 28198 173646 28250
rect 173698 28198 204158 28250
rect 204210 28198 204262 28250
rect 204314 28198 204366 28250
rect 204418 28198 218624 28250
rect 1344 28164 218624 28198
rect 1344 27466 218624 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 65918 27466
rect 65970 27414 66022 27466
rect 66074 27414 66126 27466
rect 66178 27414 96638 27466
rect 96690 27414 96742 27466
rect 96794 27414 96846 27466
rect 96898 27414 127358 27466
rect 127410 27414 127462 27466
rect 127514 27414 127566 27466
rect 127618 27414 158078 27466
rect 158130 27414 158182 27466
rect 158234 27414 158286 27466
rect 158338 27414 188798 27466
rect 188850 27414 188902 27466
rect 188954 27414 189006 27466
rect 189058 27414 218624 27466
rect 1344 27380 218624 27414
rect 1344 26682 218624 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 50558 26682
rect 50610 26630 50662 26682
rect 50714 26630 50766 26682
rect 50818 26630 81278 26682
rect 81330 26630 81382 26682
rect 81434 26630 81486 26682
rect 81538 26630 111998 26682
rect 112050 26630 112102 26682
rect 112154 26630 112206 26682
rect 112258 26630 142718 26682
rect 142770 26630 142822 26682
rect 142874 26630 142926 26682
rect 142978 26630 173438 26682
rect 173490 26630 173542 26682
rect 173594 26630 173646 26682
rect 173698 26630 204158 26682
rect 204210 26630 204262 26682
rect 204314 26630 204366 26682
rect 204418 26630 218624 26682
rect 1344 26596 218624 26630
rect 1344 25898 218624 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 65918 25898
rect 65970 25846 66022 25898
rect 66074 25846 66126 25898
rect 66178 25846 96638 25898
rect 96690 25846 96742 25898
rect 96794 25846 96846 25898
rect 96898 25846 127358 25898
rect 127410 25846 127462 25898
rect 127514 25846 127566 25898
rect 127618 25846 158078 25898
rect 158130 25846 158182 25898
rect 158234 25846 158286 25898
rect 158338 25846 188798 25898
rect 188850 25846 188902 25898
rect 188954 25846 189006 25898
rect 189058 25846 218624 25898
rect 1344 25812 218624 25846
rect 1344 25114 218624 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 50558 25114
rect 50610 25062 50662 25114
rect 50714 25062 50766 25114
rect 50818 25062 81278 25114
rect 81330 25062 81382 25114
rect 81434 25062 81486 25114
rect 81538 25062 111998 25114
rect 112050 25062 112102 25114
rect 112154 25062 112206 25114
rect 112258 25062 142718 25114
rect 142770 25062 142822 25114
rect 142874 25062 142926 25114
rect 142978 25062 173438 25114
rect 173490 25062 173542 25114
rect 173594 25062 173646 25114
rect 173698 25062 204158 25114
rect 204210 25062 204262 25114
rect 204314 25062 204366 25114
rect 204418 25062 218624 25114
rect 1344 25028 218624 25062
rect 1344 24330 218624 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 65918 24330
rect 65970 24278 66022 24330
rect 66074 24278 66126 24330
rect 66178 24278 96638 24330
rect 96690 24278 96742 24330
rect 96794 24278 96846 24330
rect 96898 24278 127358 24330
rect 127410 24278 127462 24330
rect 127514 24278 127566 24330
rect 127618 24278 158078 24330
rect 158130 24278 158182 24330
rect 158234 24278 158286 24330
rect 158338 24278 188798 24330
rect 188850 24278 188902 24330
rect 188954 24278 189006 24330
rect 189058 24278 218624 24330
rect 1344 24244 218624 24278
rect 1344 23546 218624 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 50558 23546
rect 50610 23494 50662 23546
rect 50714 23494 50766 23546
rect 50818 23494 81278 23546
rect 81330 23494 81382 23546
rect 81434 23494 81486 23546
rect 81538 23494 111998 23546
rect 112050 23494 112102 23546
rect 112154 23494 112206 23546
rect 112258 23494 142718 23546
rect 142770 23494 142822 23546
rect 142874 23494 142926 23546
rect 142978 23494 173438 23546
rect 173490 23494 173542 23546
rect 173594 23494 173646 23546
rect 173698 23494 204158 23546
rect 204210 23494 204262 23546
rect 204314 23494 204366 23546
rect 204418 23494 218624 23546
rect 1344 23460 218624 23494
rect 1344 22762 218624 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 65918 22762
rect 65970 22710 66022 22762
rect 66074 22710 66126 22762
rect 66178 22710 96638 22762
rect 96690 22710 96742 22762
rect 96794 22710 96846 22762
rect 96898 22710 127358 22762
rect 127410 22710 127462 22762
rect 127514 22710 127566 22762
rect 127618 22710 158078 22762
rect 158130 22710 158182 22762
rect 158234 22710 158286 22762
rect 158338 22710 188798 22762
rect 188850 22710 188902 22762
rect 188954 22710 189006 22762
rect 189058 22710 218624 22762
rect 1344 22676 218624 22710
rect 1344 21978 218624 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 50558 21978
rect 50610 21926 50662 21978
rect 50714 21926 50766 21978
rect 50818 21926 81278 21978
rect 81330 21926 81382 21978
rect 81434 21926 81486 21978
rect 81538 21926 111998 21978
rect 112050 21926 112102 21978
rect 112154 21926 112206 21978
rect 112258 21926 142718 21978
rect 142770 21926 142822 21978
rect 142874 21926 142926 21978
rect 142978 21926 173438 21978
rect 173490 21926 173542 21978
rect 173594 21926 173646 21978
rect 173698 21926 204158 21978
rect 204210 21926 204262 21978
rect 204314 21926 204366 21978
rect 204418 21926 218624 21978
rect 1344 21892 218624 21926
rect 1344 21194 218624 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 65918 21194
rect 65970 21142 66022 21194
rect 66074 21142 66126 21194
rect 66178 21142 96638 21194
rect 96690 21142 96742 21194
rect 96794 21142 96846 21194
rect 96898 21142 127358 21194
rect 127410 21142 127462 21194
rect 127514 21142 127566 21194
rect 127618 21142 158078 21194
rect 158130 21142 158182 21194
rect 158234 21142 158286 21194
rect 158338 21142 188798 21194
rect 188850 21142 188902 21194
rect 188954 21142 189006 21194
rect 189058 21142 218624 21194
rect 1344 21108 218624 21142
rect 1344 20410 218624 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 50558 20410
rect 50610 20358 50662 20410
rect 50714 20358 50766 20410
rect 50818 20358 81278 20410
rect 81330 20358 81382 20410
rect 81434 20358 81486 20410
rect 81538 20358 111998 20410
rect 112050 20358 112102 20410
rect 112154 20358 112206 20410
rect 112258 20358 142718 20410
rect 142770 20358 142822 20410
rect 142874 20358 142926 20410
rect 142978 20358 173438 20410
rect 173490 20358 173542 20410
rect 173594 20358 173646 20410
rect 173698 20358 204158 20410
rect 204210 20358 204262 20410
rect 204314 20358 204366 20410
rect 204418 20358 218624 20410
rect 1344 20324 218624 20358
rect 1344 19626 218624 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 65918 19626
rect 65970 19574 66022 19626
rect 66074 19574 66126 19626
rect 66178 19574 96638 19626
rect 96690 19574 96742 19626
rect 96794 19574 96846 19626
rect 96898 19574 127358 19626
rect 127410 19574 127462 19626
rect 127514 19574 127566 19626
rect 127618 19574 158078 19626
rect 158130 19574 158182 19626
rect 158234 19574 158286 19626
rect 158338 19574 188798 19626
rect 188850 19574 188902 19626
rect 188954 19574 189006 19626
rect 189058 19574 218624 19626
rect 1344 19540 218624 19574
rect 1344 18842 218624 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 50558 18842
rect 50610 18790 50662 18842
rect 50714 18790 50766 18842
rect 50818 18790 81278 18842
rect 81330 18790 81382 18842
rect 81434 18790 81486 18842
rect 81538 18790 111998 18842
rect 112050 18790 112102 18842
rect 112154 18790 112206 18842
rect 112258 18790 142718 18842
rect 142770 18790 142822 18842
rect 142874 18790 142926 18842
rect 142978 18790 173438 18842
rect 173490 18790 173542 18842
rect 173594 18790 173646 18842
rect 173698 18790 204158 18842
rect 204210 18790 204262 18842
rect 204314 18790 204366 18842
rect 204418 18790 218624 18842
rect 1344 18756 218624 18790
rect 1344 18058 218624 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 65918 18058
rect 65970 18006 66022 18058
rect 66074 18006 66126 18058
rect 66178 18006 96638 18058
rect 96690 18006 96742 18058
rect 96794 18006 96846 18058
rect 96898 18006 127358 18058
rect 127410 18006 127462 18058
rect 127514 18006 127566 18058
rect 127618 18006 158078 18058
rect 158130 18006 158182 18058
rect 158234 18006 158286 18058
rect 158338 18006 188798 18058
rect 188850 18006 188902 18058
rect 188954 18006 189006 18058
rect 189058 18006 218624 18058
rect 1344 17972 218624 18006
rect 1344 17274 218624 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 50558 17274
rect 50610 17222 50662 17274
rect 50714 17222 50766 17274
rect 50818 17222 81278 17274
rect 81330 17222 81382 17274
rect 81434 17222 81486 17274
rect 81538 17222 111998 17274
rect 112050 17222 112102 17274
rect 112154 17222 112206 17274
rect 112258 17222 142718 17274
rect 142770 17222 142822 17274
rect 142874 17222 142926 17274
rect 142978 17222 173438 17274
rect 173490 17222 173542 17274
rect 173594 17222 173646 17274
rect 173698 17222 204158 17274
rect 204210 17222 204262 17274
rect 204314 17222 204366 17274
rect 204418 17222 218624 17274
rect 1344 17188 218624 17222
rect 1344 16490 218624 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 65918 16490
rect 65970 16438 66022 16490
rect 66074 16438 66126 16490
rect 66178 16438 96638 16490
rect 96690 16438 96742 16490
rect 96794 16438 96846 16490
rect 96898 16438 127358 16490
rect 127410 16438 127462 16490
rect 127514 16438 127566 16490
rect 127618 16438 158078 16490
rect 158130 16438 158182 16490
rect 158234 16438 158286 16490
rect 158338 16438 188798 16490
rect 188850 16438 188902 16490
rect 188954 16438 189006 16490
rect 189058 16438 218624 16490
rect 1344 16404 218624 16438
rect 1344 15706 218624 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 50558 15706
rect 50610 15654 50662 15706
rect 50714 15654 50766 15706
rect 50818 15654 81278 15706
rect 81330 15654 81382 15706
rect 81434 15654 81486 15706
rect 81538 15654 111998 15706
rect 112050 15654 112102 15706
rect 112154 15654 112206 15706
rect 112258 15654 142718 15706
rect 142770 15654 142822 15706
rect 142874 15654 142926 15706
rect 142978 15654 173438 15706
rect 173490 15654 173542 15706
rect 173594 15654 173646 15706
rect 173698 15654 204158 15706
rect 204210 15654 204262 15706
rect 204314 15654 204366 15706
rect 204418 15654 218624 15706
rect 1344 15620 218624 15654
rect 1344 14922 218624 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 65918 14922
rect 65970 14870 66022 14922
rect 66074 14870 66126 14922
rect 66178 14870 96638 14922
rect 96690 14870 96742 14922
rect 96794 14870 96846 14922
rect 96898 14870 127358 14922
rect 127410 14870 127462 14922
rect 127514 14870 127566 14922
rect 127618 14870 158078 14922
rect 158130 14870 158182 14922
rect 158234 14870 158286 14922
rect 158338 14870 188798 14922
rect 188850 14870 188902 14922
rect 188954 14870 189006 14922
rect 189058 14870 218624 14922
rect 1344 14836 218624 14870
rect 1344 14138 218624 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 50558 14138
rect 50610 14086 50662 14138
rect 50714 14086 50766 14138
rect 50818 14086 81278 14138
rect 81330 14086 81382 14138
rect 81434 14086 81486 14138
rect 81538 14086 111998 14138
rect 112050 14086 112102 14138
rect 112154 14086 112206 14138
rect 112258 14086 142718 14138
rect 142770 14086 142822 14138
rect 142874 14086 142926 14138
rect 142978 14086 173438 14138
rect 173490 14086 173542 14138
rect 173594 14086 173646 14138
rect 173698 14086 204158 14138
rect 204210 14086 204262 14138
rect 204314 14086 204366 14138
rect 204418 14086 218624 14138
rect 1344 14052 218624 14086
rect 1344 13354 218624 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 65918 13354
rect 65970 13302 66022 13354
rect 66074 13302 66126 13354
rect 66178 13302 96638 13354
rect 96690 13302 96742 13354
rect 96794 13302 96846 13354
rect 96898 13302 127358 13354
rect 127410 13302 127462 13354
rect 127514 13302 127566 13354
rect 127618 13302 158078 13354
rect 158130 13302 158182 13354
rect 158234 13302 158286 13354
rect 158338 13302 188798 13354
rect 188850 13302 188902 13354
rect 188954 13302 189006 13354
rect 189058 13302 218624 13354
rect 1344 13268 218624 13302
rect 1344 12570 218624 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 50558 12570
rect 50610 12518 50662 12570
rect 50714 12518 50766 12570
rect 50818 12518 81278 12570
rect 81330 12518 81382 12570
rect 81434 12518 81486 12570
rect 81538 12518 111998 12570
rect 112050 12518 112102 12570
rect 112154 12518 112206 12570
rect 112258 12518 142718 12570
rect 142770 12518 142822 12570
rect 142874 12518 142926 12570
rect 142978 12518 173438 12570
rect 173490 12518 173542 12570
rect 173594 12518 173646 12570
rect 173698 12518 204158 12570
rect 204210 12518 204262 12570
rect 204314 12518 204366 12570
rect 204418 12518 218624 12570
rect 1344 12484 218624 12518
rect 156494 12178 156546 12190
rect 156494 12114 156546 12126
rect 163326 12066 163378 12078
rect 156034 12014 156046 12066
rect 156098 12014 156110 12066
rect 163326 12002 163378 12014
rect 1344 11786 218624 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 65918 11786
rect 65970 11734 66022 11786
rect 66074 11734 66126 11786
rect 66178 11734 96638 11786
rect 96690 11734 96742 11786
rect 96794 11734 96846 11786
rect 96898 11734 127358 11786
rect 127410 11734 127462 11786
rect 127514 11734 127566 11786
rect 127618 11734 158078 11786
rect 158130 11734 158182 11786
rect 158234 11734 158286 11786
rect 158338 11734 188798 11786
rect 188850 11734 188902 11786
rect 188954 11734 189006 11786
rect 189058 11734 218624 11786
rect 1344 11700 218624 11734
rect 156606 11618 156658 11630
rect 156606 11554 156658 11566
rect 162542 11618 162594 11630
rect 162542 11554 162594 11566
rect 146862 11506 146914 11518
rect 146862 11442 146914 11454
rect 147310 11506 147362 11518
rect 147310 11442 147362 11454
rect 149214 11506 149266 11518
rect 157726 11506 157778 11518
rect 150434 11454 150446 11506
rect 150498 11454 150510 11506
rect 155250 11454 155262 11506
rect 155314 11454 155326 11506
rect 149214 11442 149266 11454
rect 157726 11442 157778 11454
rect 164670 11506 164722 11518
rect 164670 11442 164722 11454
rect 147534 11394 147586 11406
rect 147534 11330 147586 11342
rect 148206 11394 148258 11406
rect 148206 11330 148258 11342
rect 148766 11394 148818 11406
rect 156718 11394 156770 11406
rect 155586 11342 155598 11394
rect 155650 11342 155662 11394
rect 148766 11330 148818 11342
rect 156718 11330 156770 11342
rect 157166 11394 157218 11406
rect 157166 11330 157218 11342
rect 162430 11394 162482 11406
rect 162430 11330 162482 11342
rect 163102 11394 163154 11406
rect 163102 11330 163154 11342
rect 163998 11394 164050 11406
rect 163998 11330 164050 11342
rect 150110 11282 150162 11294
rect 150110 11218 150162 11230
rect 156494 11282 156546 11294
rect 156494 11218 156546 11230
rect 163438 11282 163490 11294
rect 163438 11218 163490 11230
rect 146190 11170 146242 11182
rect 156942 11170 156994 11182
rect 147858 11118 147870 11170
rect 147922 11118 147934 11170
rect 146190 11106 146242 11118
rect 156942 11106 156994 11118
rect 162654 11170 162706 11182
rect 162654 11106 162706 11118
rect 162878 11170 162930 11182
rect 162878 11106 162930 11118
rect 163326 11170 163378 11182
rect 163326 11106 163378 11118
rect 163662 11170 163714 11182
rect 163662 11106 163714 11118
rect 163886 11170 163938 11182
rect 163886 11106 163938 11118
rect 1344 11002 218624 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 50558 11002
rect 50610 10950 50662 11002
rect 50714 10950 50766 11002
rect 50818 10950 81278 11002
rect 81330 10950 81382 11002
rect 81434 10950 81486 11002
rect 81538 10950 111998 11002
rect 112050 10950 112102 11002
rect 112154 10950 112206 11002
rect 112258 10950 142718 11002
rect 142770 10950 142822 11002
rect 142874 10950 142926 11002
rect 142978 10950 173438 11002
rect 173490 10950 173542 11002
rect 173594 10950 173646 11002
rect 173698 10950 204158 11002
rect 204210 10950 204262 11002
rect 204314 10950 204366 11002
rect 204418 10950 218624 11002
rect 1344 10916 218624 10950
rect 147870 10834 147922 10846
rect 147870 10770 147922 10782
rect 161534 10834 161586 10846
rect 161534 10770 161586 10782
rect 162318 10834 162370 10846
rect 162318 10770 162370 10782
rect 162990 10834 163042 10846
rect 162990 10770 163042 10782
rect 163550 10834 163602 10846
rect 163550 10770 163602 10782
rect 163774 10834 163826 10846
rect 163774 10770 163826 10782
rect 164446 10834 164498 10846
rect 164446 10770 164498 10782
rect 160526 10722 160578 10734
rect 154914 10670 154926 10722
rect 154978 10670 154990 10722
rect 156146 10670 156158 10722
rect 156210 10670 156222 10722
rect 160526 10658 160578 10670
rect 160750 10722 160802 10734
rect 160750 10658 160802 10670
rect 162094 10722 162146 10734
rect 162094 10658 162146 10670
rect 163998 10722 164050 10734
rect 163998 10658 164050 10670
rect 148206 10610 148258 10622
rect 149662 10610 149714 10622
rect 149202 10558 149214 10610
rect 149266 10558 149278 10610
rect 148206 10546 148258 10558
rect 149662 10546 149714 10558
rect 151230 10610 151282 10622
rect 151230 10546 151282 10558
rect 153134 10610 153186 10622
rect 160078 10610 160130 10622
rect 155698 10558 155710 10610
rect 155762 10558 155774 10610
rect 156034 10558 156046 10610
rect 156098 10558 156110 10610
rect 153134 10546 153186 10558
rect 160078 10546 160130 10558
rect 160302 10610 160354 10622
rect 160302 10546 160354 10558
rect 161198 10610 161250 10622
rect 161198 10546 161250 10558
rect 161982 10610 162034 10622
rect 161982 10546 162034 10558
rect 162542 10610 162594 10622
rect 162542 10546 162594 10558
rect 163326 10610 163378 10622
rect 163326 10546 163378 10558
rect 147534 10498 147586 10510
rect 147534 10434 147586 10446
rect 148766 10498 148818 10510
rect 148766 10434 148818 10446
rect 151790 10498 151842 10510
rect 162654 10498 162706 10510
rect 153570 10446 153582 10498
rect 153634 10446 153646 10498
rect 154578 10446 154590 10498
rect 154642 10446 154654 10498
rect 151790 10434 151842 10446
rect 162654 10434 162706 10446
rect 160190 10386 160242 10398
rect 160190 10322 160242 10334
rect 163438 10386 163490 10398
rect 163438 10322 163490 10334
rect 1344 10218 218624 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 65918 10218
rect 65970 10166 66022 10218
rect 66074 10166 66126 10218
rect 66178 10166 96638 10218
rect 96690 10166 96742 10218
rect 96794 10166 96846 10218
rect 96898 10166 127358 10218
rect 127410 10166 127462 10218
rect 127514 10166 127566 10218
rect 127618 10166 158078 10218
rect 158130 10166 158182 10218
rect 158234 10166 158286 10218
rect 158338 10166 188798 10218
rect 188850 10166 188902 10218
rect 188954 10166 189006 10218
rect 189058 10166 218624 10218
rect 1344 10132 218624 10166
rect 139794 9998 139806 10050
rect 139858 10047 139870 10050
rect 140354 10047 140366 10050
rect 139858 10001 140366 10047
rect 139858 9998 139870 10001
rect 140354 9998 140366 10001
rect 140418 9998 140430 10050
rect 139134 9938 139186 9950
rect 139134 9874 139186 9886
rect 139806 9938 139858 9950
rect 139806 9874 139858 9886
rect 140366 9938 140418 9950
rect 140366 9874 140418 9886
rect 148206 9938 148258 9950
rect 148206 9874 148258 9886
rect 157950 9938 158002 9950
rect 157950 9874 158002 9886
rect 161086 9938 161138 9950
rect 161086 9874 161138 9886
rect 140702 9826 140754 9838
rect 140702 9762 140754 9774
rect 148542 9826 148594 9838
rect 148542 9762 148594 9774
rect 149774 9826 149826 9838
rect 151902 9826 151954 9838
rect 151554 9774 151566 9826
rect 151618 9774 151630 9826
rect 149774 9762 149826 9774
rect 151902 9762 151954 9774
rect 152462 9826 152514 9838
rect 152462 9762 152514 9774
rect 154814 9826 154866 9838
rect 154814 9762 154866 9774
rect 155598 9826 155650 9838
rect 155598 9762 155650 9774
rect 155934 9826 155986 9838
rect 155934 9762 155986 9774
rect 156158 9826 156210 9838
rect 156158 9762 156210 9774
rect 156830 9826 156882 9838
rect 156830 9762 156882 9774
rect 157502 9826 157554 9838
rect 157502 9762 157554 9774
rect 150558 9714 150610 9726
rect 150558 9650 150610 9662
rect 155150 9714 155202 9726
rect 155150 9650 155202 9662
rect 157054 9714 157106 9726
rect 157054 9650 157106 9662
rect 161534 9714 161586 9726
rect 161534 9650 161586 9662
rect 161870 9714 161922 9726
rect 161870 9650 161922 9662
rect 141486 9602 141538 9614
rect 141486 9538 141538 9550
rect 148654 9602 148706 9614
rect 148654 9538 148706 9550
rect 149998 9602 150050 9614
rect 149998 9538 150050 9550
rect 154030 9602 154082 9614
rect 154030 9538 154082 9550
rect 155710 9602 155762 9614
rect 155710 9538 155762 9550
rect 156270 9602 156322 9614
rect 156270 9538 156322 9550
rect 156718 9602 156770 9614
rect 156718 9538 156770 9550
rect 157278 9602 157330 9614
rect 157278 9538 157330 9550
rect 1344 9434 218624 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 50558 9434
rect 50610 9382 50662 9434
rect 50714 9382 50766 9434
rect 50818 9382 81278 9434
rect 81330 9382 81382 9434
rect 81434 9382 81486 9434
rect 81538 9382 111998 9434
rect 112050 9382 112102 9434
rect 112154 9382 112206 9434
rect 112258 9382 142718 9434
rect 142770 9382 142822 9434
rect 142874 9382 142926 9434
rect 142978 9382 173438 9434
rect 173490 9382 173542 9434
rect 173594 9382 173646 9434
rect 173698 9382 204158 9434
rect 204210 9382 204262 9434
rect 204314 9382 204366 9434
rect 204418 9382 218624 9434
rect 1344 9348 218624 9382
rect 138686 9266 138738 9278
rect 138686 9202 138738 9214
rect 139582 9266 139634 9278
rect 139582 9202 139634 9214
rect 148430 9266 148482 9278
rect 148430 9202 148482 9214
rect 150110 9266 150162 9278
rect 150110 9202 150162 9214
rect 151566 9266 151618 9278
rect 151566 9202 151618 9214
rect 156046 9266 156098 9278
rect 156046 9202 156098 9214
rect 157166 9266 157218 9278
rect 157166 9202 157218 9214
rect 135326 9154 135378 9166
rect 148542 9154 148594 9166
rect 135986 9102 135998 9154
rect 136050 9102 136062 9154
rect 138226 9102 138238 9154
rect 138290 9102 138302 9154
rect 140242 9102 140254 9154
rect 140306 9102 140318 9154
rect 140914 9102 140926 9154
rect 140978 9102 140990 9154
rect 135326 9090 135378 9102
rect 148542 9090 148594 9102
rect 151006 9154 151058 9166
rect 151006 9090 151058 9102
rect 153358 9154 153410 9166
rect 153358 9090 153410 9102
rect 134542 9042 134594 9054
rect 149326 9042 149378 9054
rect 150670 9042 150722 9054
rect 135538 8990 135550 9042
rect 135602 8990 135614 9042
rect 137666 8990 137678 9042
rect 137730 8990 137742 9042
rect 140802 8990 140814 9042
rect 140866 8990 140878 9042
rect 149538 8990 149550 9042
rect 149602 8990 149614 9042
rect 134542 8978 134594 8990
rect 149326 8978 149378 8990
rect 150670 8978 150722 8990
rect 152126 9042 152178 9054
rect 153906 8990 153918 9042
rect 153970 8990 153982 9042
rect 152126 8978 152178 8990
rect 149662 8930 149714 8942
rect 139122 8878 139134 8930
rect 139186 8878 139198 8930
rect 156482 8878 156494 8930
rect 156546 8878 156558 8930
rect 149662 8866 149714 8878
rect 1344 8650 218624 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 65918 8650
rect 65970 8598 66022 8650
rect 66074 8598 66126 8650
rect 66178 8598 96638 8650
rect 96690 8598 96742 8650
rect 96794 8598 96846 8650
rect 96898 8598 127358 8650
rect 127410 8598 127462 8650
rect 127514 8598 127566 8650
rect 127618 8598 158078 8650
rect 158130 8598 158182 8650
rect 158234 8598 158286 8650
rect 158338 8598 188798 8650
rect 188850 8598 188902 8650
rect 188954 8598 189006 8650
rect 189058 8598 218624 8650
rect 1344 8564 218624 8598
rect 153010 8430 153022 8482
rect 153074 8479 153086 8482
rect 153074 8433 153519 8479
rect 153074 8430 153086 8433
rect 132862 8370 132914 8382
rect 147870 8370 147922 8382
rect 144722 8318 144734 8370
rect 144786 8318 144798 8370
rect 132862 8306 132914 8318
rect 147870 8306 147922 8318
rect 148542 8370 148594 8382
rect 148542 8306 148594 8318
rect 148766 8370 148818 8382
rect 148766 8306 148818 8318
rect 149886 8370 149938 8382
rect 149886 8306 149938 8318
rect 152798 8370 152850 8382
rect 153473 8367 153519 8433
rect 153694 8370 153746 8382
rect 153570 8367 153582 8370
rect 153473 8321 153582 8367
rect 153570 8318 153582 8321
rect 153634 8318 153646 8370
rect 152798 8306 152850 8318
rect 153694 8306 153746 8318
rect 150222 8258 150274 8270
rect 133074 8206 133086 8258
rect 133138 8206 133150 8258
rect 135538 8206 135550 8258
rect 135602 8206 135614 8258
rect 139458 8206 139470 8258
rect 139522 8206 139534 8258
rect 140914 8206 140926 8258
rect 140978 8206 140990 8258
rect 150222 8194 150274 8206
rect 152350 8258 152402 8270
rect 152350 8194 152402 8206
rect 162430 8258 162482 8270
rect 162430 8194 162482 8206
rect 150670 8146 150722 8158
rect 133186 8094 133198 8146
rect 133250 8094 133262 8146
rect 135762 8094 135774 8146
rect 135826 8094 135838 8146
rect 139570 8094 139582 8146
rect 139634 8094 139646 8146
rect 142146 8094 142158 8146
rect 142210 8094 142222 8146
rect 150670 8082 150722 8094
rect 136334 8034 136386 8046
rect 136334 7970 136386 7982
rect 138462 8034 138514 8046
rect 143278 8034 143330 8046
rect 140130 7982 140142 8034
rect 140194 7982 140206 8034
rect 138462 7970 138514 7982
rect 143278 7970 143330 7982
rect 144062 8034 144114 8046
rect 144062 7970 144114 7982
rect 145182 8034 145234 8046
rect 150222 8034 150274 8046
rect 153358 8034 153410 8046
rect 148194 7982 148206 8034
rect 148258 7982 148270 8034
rect 152002 7982 152014 8034
rect 152066 7982 152078 8034
rect 145182 7970 145234 7982
rect 150222 7970 150274 7982
rect 153358 7970 153410 7982
rect 154702 8034 154754 8046
rect 162754 7982 162766 8034
rect 162818 7982 162830 8034
rect 154702 7970 154754 7982
rect 1344 7866 218624 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 50558 7866
rect 50610 7814 50662 7866
rect 50714 7814 50766 7866
rect 50818 7814 81278 7866
rect 81330 7814 81382 7866
rect 81434 7814 81486 7866
rect 81538 7814 111998 7866
rect 112050 7814 112102 7866
rect 112154 7814 112206 7866
rect 112258 7814 142718 7866
rect 142770 7814 142822 7866
rect 142874 7814 142926 7866
rect 142978 7814 173438 7866
rect 173490 7814 173542 7866
rect 173594 7814 173646 7866
rect 173698 7814 204158 7866
rect 204210 7814 204262 7866
rect 204314 7814 204366 7866
rect 204418 7814 218624 7866
rect 1344 7780 218624 7814
rect 151902 7698 151954 7710
rect 132738 7646 132750 7698
rect 132802 7646 132814 7698
rect 136210 7646 136222 7698
rect 136274 7646 136286 7698
rect 140018 7646 140030 7698
rect 140082 7646 140094 7698
rect 147858 7646 147870 7698
rect 147922 7646 147934 7698
rect 151902 7634 151954 7646
rect 153134 7698 153186 7710
rect 153134 7634 153186 7646
rect 153806 7698 153858 7710
rect 153806 7634 153858 7646
rect 160638 7698 160690 7710
rect 160638 7634 160690 7646
rect 151342 7586 151394 7598
rect 132514 7534 132526 7586
rect 132578 7534 132590 7586
rect 133970 7534 133982 7586
rect 134034 7534 134046 7586
rect 135650 7534 135662 7586
rect 135714 7534 135726 7586
rect 138226 7534 138238 7586
rect 138290 7534 138302 7586
rect 139458 7534 139470 7586
rect 139522 7534 139534 7586
rect 142930 7534 142942 7586
rect 142994 7534 143006 7586
rect 148082 7534 148094 7586
rect 148146 7534 148158 7586
rect 151342 7522 151394 7534
rect 151678 7586 151730 7598
rect 151678 7522 151730 7534
rect 152686 7586 152738 7598
rect 152686 7522 152738 7534
rect 161758 7586 161810 7598
rect 161758 7522 161810 7534
rect 162766 7586 162818 7598
rect 162766 7522 162818 7534
rect 163550 7586 163602 7598
rect 163550 7522 163602 7534
rect 141822 7474 141874 7486
rect 150782 7474 150834 7486
rect 131730 7422 131742 7474
rect 131794 7422 131806 7474
rect 134194 7422 134206 7474
rect 134258 7422 134270 7474
rect 135538 7422 135550 7474
rect 135602 7422 135614 7474
rect 137666 7422 137678 7474
rect 137730 7422 137742 7474
rect 139122 7422 139134 7474
rect 139186 7422 139198 7474
rect 140578 7422 140590 7474
rect 140642 7422 140654 7474
rect 144050 7422 144062 7474
rect 144114 7422 144126 7474
rect 145730 7422 145742 7474
rect 145794 7422 145806 7474
rect 146066 7422 146078 7474
rect 146130 7422 146142 7474
rect 146402 7422 146414 7474
rect 146466 7422 146478 7474
rect 147634 7422 147646 7474
rect 147698 7422 147710 7474
rect 149314 7422 149326 7474
rect 149378 7422 149390 7474
rect 141822 7410 141874 7422
rect 150782 7410 150834 7422
rect 150894 7474 150946 7486
rect 150894 7410 150946 7422
rect 151118 7474 151170 7486
rect 151118 7410 151170 7422
rect 152126 7474 152178 7486
rect 152126 7410 152178 7422
rect 152350 7474 152402 7486
rect 152350 7410 152402 7422
rect 152910 7474 152962 7486
rect 152910 7410 152962 7422
rect 153246 7474 153298 7486
rect 153246 7410 153298 7422
rect 161422 7474 161474 7486
rect 161422 7410 161474 7422
rect 162206 7474 162258 7486
rect 162990 7474 163042 7486
rect 162530 7422 162542 7474
rect 162594 7422 162606 7474
rect 163314 7422 163326 7474
rect 163378 7422 163390 7474
rect 162206 7410 162258 7422
rect 162990 7410 163042 7422
rect 150110 7362 150162 7374
rect 150110 7298 150162 7310
rect 151454 7362 151506 7374
rect 151454 7298 151506 7310
rect 152462 7362 152514 7374
rect 152462 7298 152514 7310
rect 154254 7362 154306 7374
rect 154254 7298 154306 7310
rect 154814 7362 154866 7374
rect 154814 7298 154866 7310
rect 155150 7362 155202 7374
rect 155150 7298 155202 7310
rect 161086 7362 161138 7374
rect 161086 7298 161138 7310
rect 164110 7362 164162 7374
rect 164110 7298 164162 7310
rect 152798 7250 152850 7262
rect 152798 7186 152850 7198
rect 162878 7250 162930 7262
rect 162878 7186 162930 7198
rect 163662 7250 163714 7262
rect 163662 7186 163714 7198
rect 1344 7082 218624 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 65918 7082
rect 65970 7030 66022 7082
rect 66074 7030 66126 7082
rect 66178 7030 96638 7082
rect 96690 7030 96742 7082
rect 96794 7030 96846 7082
rect 96898 7030 127358 7082
rect 127410 7030 127462 7082
rect 127514 7030 127566 7082
rect 127618 7030 158078 7082
rect 158130 7030 158182 7082
rect 158234 7030 158286 7082
rect 158338 7030 188798 7082
rect 188850 7030 188902 7082
rect 188954 7030 189006 7082
rect 189058 7030 218624 7082
rect 1344 6996 218624 7030
rect 151902 6802 151954 6814
rect 161534 6802 161586 6814
rect 155362 6750 155374 6802
rect 155426 6750 155438 6802
rect 160626 6750 160638 6802
rect 160690 6750 160702 6802
rect 151902 6738 151954 6750
rect 161534 6738 161586 6750
rect 162766 6802 162818 6814
rect 162766 6738 162818 6750
rect 137230 6690 137282 6702
rect 133074 6638 133086 6690
rect 133138 6638 133150 6690
rect 135202 6638 135214 6690
rect 135266 6638 135278 6690
rect 136322 6638 136334 6690
rect 136386 6638 136398 6690
rect 137230 6626 137282 6638
rect 138238 6690 138290 6702
rect 145406 6690 145458 6702
rect 139010 6638 139022 6690
rect 139074 6638 139086 6690
rect 141810 6638 141822 6690
rect 141874 6638 141886 6690
rect 142482 6638 142494 6690
rect 142546 6638 142558 6690
rect 142930 6638 142942 6690
rect 142994 6638 143006 6690
rect 138238 6626 138290 6638
rect 145406 6626 145458 6638
rect 145854 6690 145906 6702
rect 145854 6626 145906 6638
rect 147646 6690 147698 6702
rect 147646 6626 147698 6638
rect 147982 6690 148034 6702
rect 160974 6690 161026 6702
rect 148642 6638 148654 6690
rect 148706 6638 148718 6690
rect 149986 6638 149998 6690
rect 150050 6638 150062 6690
rect 150322 6638 150334 6690
rect 150386 6638 150398 6690
rect 151106 6638 151118 6690
rect 151170 6638 151182 6690
rect 153346 6638 153358 6690
rect 153410 6638 153422 6690
rect 155586 6638 155598 6690
rect 155650 6638 155662 6690
rect 155810 6638 155822 6690
rect 155874 6638 155886 6690
rect 147982 6626 148034 6638
rect 160974 6626 161026 6638
rect 162654 6690 162706 6702
rect 162654 6626 162706 6638
rect 163886 6690 163938 6702
rect 163886 6626 163938 6638
rect 164334 6690 164386 6702
rect 164334 6626 164386 6638
rect 144622 6578 144674 6590
rect 160302 6578 160354 6590
rect 133186 6526 133198 6578
rect 133250 6526 133262 6578
rect 135762 6526 135774 6578
rect 135826 6526 135838 6578
rect 140354 6526 140366 6578
rect 140418 6526 140430 6578
rect 140690 6526 140702 6578
rect 140754 6526 140766 6578
rect 152114 6526 152126 6578
rect 152178 6526 152190 6578
rect 156594 6526 156606 6578
rect 156658 6526 156670 6578
rect 144622 6514 144674 6526
rect 160302 6514 160354 6526
rect 161422 6578 161474 6590
rect 161422 6514 161474 6526
rect 162878 6578 162930 6590
rect 162878 6514 162930 6526
rect 137902 6466 137954 6478
rect 144286 6466 144338 6478
rect 134642 6414 134654 6466
rect 134706 6414 134718 6466
rect 138898 6414 138910 6466
rect 138962 6414 138974 6466
rect 137902 6402 137954 6414
rect 144286 6402 144338 6414
rect 147310 6466 147362 6478
rect 154030 6466 154082 6478
rect 148306 6414 148318 6466
rect 148370 6414 148382 6466
rect 147310 6402 147362 6414
rect 154030 6402 154082 6414
rect 159966 6466 160018 6478
rect 159966 6402 160018 6414
rect 160526 6466 160578 6478
rect 160526 6402 160578 6414
rect 160750 6466 160802 6478
rect 160750 6402 160802 6414
rect 161646 6466 161698 6478
rect 161646 6402 161698 6414
rect 163102 6466 163154 6478
rect 163102 6402 163154 6414
rect 163774 6466 163826 6478
rect 163774 6402 163826 6414
rect 164446 6466 164498 6478
rect 164446 6402 164498 6414
rect 164558 6466 164610 6478
rect 164558 6402 164610 6414
rect 165118 6466 165170 6478
rect 165118 6402 165170 6414
rect 1344 6298 218624 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 50558 6298
rect 50610 6246 50662 6298
rect 50714 6246 50766 6298
rect 50818 6246 81278 6298
rect 81330 6246 81382 6298
rect 81434 6246 81486 6298
rect 81538 6246 111998 6298
rect 112050 6246 112102 6298
rect 112154 6246 112206 6298
rect 112258 6246 142718 6298
rect 142770 6246 142822 6298
rect 142874 6246 142926 6298
rect 142978 6246 173438 6298
rect 173490 6246 173542 6298
rect 173594 6246 173646 6298
rect 173698 6246 204158 6298
rect 204210 6246 204262 6298
rect 204314 6246 204366 6298
rect 204418 6246 218624 6298
rect 1344 6212 218624 6246
rect 135550 6130 135602 6142
rect 149662 6130 149714 6142
rect 138002 6078 138014 6130
rect 138066 6078 138078 6130
rect 145282 6078 145294 6130
rect 145346 6078 145358 6130
rect 135550 6066 135602 6078
rect 149662 6066 149714 6078
rect 156830 6130 156882 6142
rect 156830 6066 156882 6078
rect 157950 6130 158002 6142
rect 157950 6066 158002 6078
rect 159294 6130 159346 6142
rect 159854 6130 159906 6142
rect 159618 6078 159630 6130
rect 159682 6078 159694 6130
rect 159294 6066 159346 6078
rect 159854 6066 159906 6078
rect 161198 6130 161250 6142
rect 161198 6066 161250 6078
rect 162318 6130 162370 6142
rect 162318 6066 162370 6078
rect 164894 6130 164946 6142
rect 164894 6066 164946 6078
rect 149886 6018 149938 6030
rect 137218 5966 137230 6018
rect 137282 5966 137294 6018
rect 139794 5966 139806 6018
rect 139858 5966 139870 6018
rect 145058 5966 145070 6018
rect 145122 5966 145134 6018
rect 149886 5954 149938 5966
rect 151454 6018 151506 6030
rect 160638 6018 160690 6030
rect 152674 5966 152686 6018
rect 152738 5966 152750 6018
rect 154690 5966 154702 6018
rect 154754 5966 154766 6018
rect 160402 5966 160414 6018
rect 160466 5966 160478 6018
rect 151454 5954 151506 5966
rect 160638 5954 160690 5966
rect 162990 6018 163042 6030
rect 163998 6018 164050 6030
rect 163202 5966 163214 6018
rect 163266 5966 163278 6018
rect 162990 5954 163042 5966
rect 163998 5954 164050 5966
rect 139134 5906 139186 5918
rect 141822 5906 141874 5918
rect 149438 5906 149490 5918
rect 136434 5854 136446 5906
rect 136498 5854 136510 5906
rect 138898 5854 138910 5906
rect 138962 5854 138974 5906
rect 140130 5854 140142 5906
rect 140194 5854 140206 5906
rect 143938 5854 143950 5906
rect 144002 5854 144014 5906
rect 146066 5854 146078 5906
rect 146130 5854 146142 5906
rect 146738 5854 146750 5906
rect 146802 5854 146814 5906
rect 147186 5854 147198 5906
rect 147250 5854 147262 5906
rect 148530 5854 148542 5906
rect 148594 5854 148606 5906
rect 139134 5842 139186 5854
rect 141822 5842 141874 5854
rect 149438 5842 149490 5854
rect 150110 5906 150162 5918
rect 160750 5906 160802 5918
rect 151330 5854 151342 5906
rect 151394 5854 151406 5906
rect 152114 5854 152126 5906
rect 152178 5854 152190 5906
rect 152450 5854 152462 5906
rect 152514 5854 152526 5906
rect 153906 5854 153918 5906
rect 153970 5854 153982 5906
rect 154130 5854 154142 5906
rect 154194 5854 154206 5906
rect 156370 5854 156382 5906
rect 156434 5854 156446 5906
rect 160178 5854 160190 5906
rect 160242 5854 160254 5906
rect 150110 5842 150162 5854
rect 160750 5842 160802 5854
rect 161758 5906 161810 5918
rect 161758 5842 161810 5854
rect 162542 5906 162594 5918
rect 162542 5842 162594 5854
rect 163326 5906 163378 5918
rect 163326 5842 163378 5854
rect 163550 5906 163602 5918
rect 163550 5842 163602 5854
rect 164110 5906 164162 5918
rect 164110 5842 164162 5854
rect 164222 5906 164274 5918
rect 164222 5842 164274 5854
rect 164446 5906 164498 5918
rect 164446 5842 164498 5854
rect 165118 5906 165170 5918
rect 165118 5842 165170 5854
rect 165566 5906 165618 5918
rect 165566 5842 165618 5854
rect 135102 5794 135154 5806
rect 140590 5794 140642 5806
rect 149102 5794 149154 5806
rect 139458 5742 139470 5794
rect 139522 5742 139534 5794
rect 141250 5742 141262 5794
rect 141314 5742 141326 5794
rect 135102 5730 135154 5742
rect 140590 5730 140642 5742
rect 149102 5730 149154 5742
rect 150222 5794 150274 5806
rect 150222 5730 150274 5742
rect 150782 5794 150834 5806
rect 150782 5730 150834 5742
rect 155934 5794 155986 5806
rect 155934 5730 155986 5742
rect 157390 5794 157442 5806
rect 157390 5730 157442 5742
rect 165006 5794 165058 5806
rect 165006 5730 165058 5742
rect 153122 5630 153134 5682
rect 153186 5630 153198 5682
rect 1344 5514 218624 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 65918 5514
rect 65970 5462 66022 5514
rect 66074 5462 66126 5514
rect 66178 5462 96638 5514
rect 96690 5462 96742 5514
rect 96794 5462 96846 5514
rect 96898 5462 127358 5514
rect 127410 5462 127462 5514
rect 127514 5462 127566 5514
rect 127618 5462 158078 5514
rect 158130 5462 158182 5514
rect 158234 5462 158286 5514
rect 158338 5462 188798 5514
rect 188850 5462 188902 5514
rect 188954 5462 189006 5514
rect 189058 5462 218624 5514
rect 1344 5428 218624 5462
rect 130510 5346 130562 5358
rect 130510 5282 130562 5294
rect 131294 5346 131346 5358
rect 131294 5282 131346 5294
rect 131742 5346 131794 5358
rect 131742 5282 131794 5294
rect 133758 5346 133810 5358
rect 133758 5282 133810 5294
rect 134206 5346 134258 5358
rect 134206 5282 134258 5294
rect 134542 5346 134594 5358
rect 134542 5282 134594 5294
rect 135774 5346 135826 5358
rect 135774 5282 135826 5294
rect 152574 5346 152626 5358
rect 152574 5282 152626 5294
rect 153022 5346 153074 5358
rect 153022 5282 153074 5294
rect 155150 5346 155202 5358
rect 155150 5282 155202 5294
rect 156382 5346 156434 5358
rect 156382 5282 156434 5294
rect 6414 5234 6466 5246
rect 6414 5170 6466 5182
rect 49758 5234 49810 5246
rect 49758 5170 49810 5182
rect 52110 5234 52162 5246
rect 52110 5170 52162 5182
rect 55134 5234 55186 5246
rect 55134 5170 55186 5182
rect 57822 5234 57874 5246
rect 57822 5170 57874 5182
rect 59950 5234 60002 5246
rect 59950 5170 60002 5182
rect 63198 5234 63250 5246
rect 63198 5170 63250 5182
rect 65886 5234 65938 5246
rect 65886 5170 65938 5182
rect 68574 5234 68626 5246
rect 68574 5170 68626 5182
rect 92766 5234 92818 5246
rect 92766 5170 92818 5182
rect 93774 5234 93826 5246
rect 98366 5234 98418 5246
rect 97458 5182 97470 5234
rect 97522 5182 97534 5234
rect 93774 5170 93826 5182
rect 98366 5170 98418 5182
rect 102062 5234 102114 5246
rect 102062 5170 102114 5182
rect 105534 5234 105586 5246
rect 105534 5170 105586 5182
rect 106542 5234 106594 5246
rect 110798 5234 110850 5246
rect 109218 5182 109230 5234
rect 109282 5182 109294 5234
rect 110338 5182 110350 5234
rect 110402 5182 110414 5234
rect 106542 5170 106594 5182
rect 110798 5170 110850 5182
rect 113374 5234 113426 5246
rect 113374 5170 113426 5182
rect 114382 5234 114434 5246
rect 118526 5234 118578 5246
rect 117618 5182 117630 5234
rect 117682 5182 117694 5234
rect 114382 5170 114434 5182
rect 118526 5170 118578 5182
rect 121214 5234 121266 5246
rect 121214 5170 121266 5182
rect 122222 5234 122274 5246
rect 122222 5170 122274 5182
rect 125582 5234 125634 5246
rect 125582 5170 125634 5182
rect 126590 5234 126642 5246
rect 126590 5170 126642 5182
rect 130062 5234 130114 5246
rect 130062 5170 130114 5182
rect 130398 5234 130450 5246
rect 130398 5170 130450 5182
rect 132078 5234 132130 5246
rect 132078 5170 132130 5182
rect 132638 5234 132690 5246
rect 132638 5170 132690 5182
rect 133422 5234 133474 5246
rect 145406 5234 145458 5246
rect 137442 5182 137454 5234
rect 137506 5182 137518 5234
rect 133422 5170 133474 5182
rect 145406 5170 145458 5182
rect 145854 5234 145906 5246
rect 145854 5170 145906 5182
rect 157950 5234 158002 5246
rect 157950 5170 158002 5182
rect 161870 5234 161922 5246
rect 161870 5170 161922 5182
rect 162878 5234 162930 5246
rect 162878 5170 162930 5182
rect 5966 5122 6018 5134
rect 5966 5058 6018 5070
rect 50094 5122 50146 5134
rect 50094 5058 50146 5070
rect 52782 5122 52834 5134
rect 52782 5058 52834 5070
rect 55470 5122 55522 5134
rect 55470 5058 55522 5070
rect 58158 5122 58210 5134
rect 58158 5058 58210 5070
rect 60846 5122 60898 5134
rect 60846 5058 60898 5070
rect 63534 5122 63586 5134
rect 63534 5058 63586 5070
rect 66222 5122 66274 5134
rect 66222 5058 66274 5070
rect 68910 5122 68962 5134
rect 68910 5058 68962 5070
rect 93326 5122 93378 5134
rect 93326 5058 93378 5070
rect 97918 5122 97970 5134
rect 97918 5058 97970 5070
rect 101614 5122 101666 5134
rect 101614 5058 101666 5070
rect 106094 5122 106146 5134
rect 106094 5058 106146 5070
rect 109678 5122 109730 5134
rect 109678 5058 109730 5070
rect 110014 5122 110066 5134
rect 110014 5058 110066 5070
rect 113934 5122 113986 5134
rect 113934 5058 113986 5070
rect 118078 5122 118130 5134
rect 118078 5058 118130 5070
rect 121774 5122 121826 5134
rect 121774 5058 121826 5070
rect 126142 5122 126194 5134
rect 126142 5058 126194 5070
rect 131182 5122 131234 5134
rect 131182 5058 131234 5070
rect 133646 5122 133698 5134
rect 133646 5058 133698 5070
rect 135326 5122 135378 5134
rect 144958 5122 145010 5134
rect 152014 5122 152066 5134
rect 136882 5070 136894 5122
rect 136946 5070 136958 5122
rect 138114 5070 138126 5122
rect 138178 5070 138190 5122
rect 138898 5070 138910 5122
rect 138962 5070 138974 5122
rect 141810 5070 141822 5122
rect 141874 5070 141886 5122
rect 142482 5070 142494 5122
rect 142546 5070 142558 5122
rect 143042 5070 143054 5122
rect 143106 5070 143118 5122
rect 144274 5070 144286 5122
rect 144338 5070 144350 5122
rect 146738 5070 146750 5122
rect 146802 5070 146814 5122
rect 148978 5070 148990 5122
rect 149042 5070 149054 5122
rect 150322 5070 150334 5122
rect 150386 5070 150398 5122
rect 150546 5070 150558 5122
rect 150610 5070 150622 5122
rect 135326 5058 135378 5070
rect 144958 5058 145010 5070
rect 152014 5058 152066 5070
rect 152238 5122 152290 5134
rect 152238 5058 152290 5070
rect 152574 5122 152626 5134
rect 153694 5122 153746 5134
rect 153458 5070 153470 5122
rect 153522 5070 153534 5122
rect 152574 5058 152626 5070
rect 153694 5058 153746 5070
rect 154030 5122 154082 5134
rect 155374 5122 155426 5134
rect 154578 5070 154590 5122
rect 154642 5070 154654 5122
rect 154030 5058 154082 5070
rect 155374 5058 155426 5070
rect 155598 5122 155650 5134
rect 155598 5058 155650 5070
rect 155710 5122 155762 5134
rect 155710 5058 155762 5070
rect 156158 5122 156210 5134
rect 156158 5058 156210 5070
rect 156718 5122 156770 5134
rect 156718 5058 156770 5070
rect 157166 5122 157218 5134
rect 157166 5058 157218 5070
rect 157278 5122 157330 5134
rect 157278 5058 157330 5070
rect 157390 5122 157442 5134
rect 161086 5122 161138 5134
rect 157826 5070 157838 5122
rect 157890 5070 157902 5122
rect 160514 5070 160526 5122
rect 160578 5070 160590 5122
rect 157390 5058 157442 5070
rect 161086 5058 161138 5070
rect 161534 5122 161586 5134
rect 161534 5058 161586 5070
rect 162318 5122 162370 5134
rect 162318 5058 162370 5070
rect 162766 5122 162818 5134
rect 162766 5058 162818 5070
rect 163326 5122 163378 5134
rect 163326 5058 163378 5070
rect 163662 5122 163714 5134
rect 163662 5058 163714 5070
rect 163774 5122 163826 5134
rect 163774 5058 163826 5070
rect 163998 5122 164050 5134
rect 163998 5058 164050 5070
rect 164782 5122 164834 5134
rect 164782 5058 164834 5070
rect 165230 5122 165282 5134
rect 165230 5058 165282 5070
rect 165678 5122 165730 5134
rect 165678 5058 165730 5070
rect 166126 5122 166178 5134
rect 166126 5058 166178 5070
rect 166238 5122 166290 5134
rect 166238 5058 166290 5070
rect 101054 5010 101106 5022
rect 101054 4946 101106 4958
rect 131630 5010 131682 5022
rect 131630 4946 131682 4958
rect 132190 5010 132242 5022
rect 132190 4946 132242 4958
rect 134094 5010 134146 5022
rect 134094 4946 134146 4958
rect 135662 5010 135714 5022
rect 152462 5010 152514 5022
rect 158286 5010 158338 5022
rect 162990 5010 163042 5022
rect 136994 4958 137006 5010
rect 137058 4958 137070 5010
rect 138002 4958 138014 5010
rect 138066 4958 138078 5010
rect 140354 4958 140366 5010
rect 140418 4958 140430 5010
rect 140690 4958 140702 5010
rect 140754 4958 140766 5010
rect 148194 4958 148206 5010
rect 148258 4958 148270 5010
rect 148530 4958 148542 5010
rect 148594 4958 148606 5010
rect 153906 4958 153918 5010
rect 153970 4958 153982 5010
rect 160290 4958 160302 5010
rect 160354 4958 160366 5010
rect 161746 4958 161758 5010
rect 161810 4958 161822 5010
rect 135662 4946 135714 4958
rect 152462 4946 152514 4958
rect 158286 4946 158338 4958
rect 162990 4946 163042 4958
rect 5630 4898 5682 4910
rect 5630 4834 5682 4846
rect 50430 4898 50482 4910
rect 50430 4834 50482 4846
rect 53118 4898 53170 4910
rect 53118 4834 53170 4846
rect 55806 4898 55858 4910
rect 55806 4834 55858 4846
rect 58494 4898 58546 4910
rect 58494 4834 58546 4846
rect 61182 4898 61234 4910
rect 61182 4834 61234 4846
rect 63870 4898 63922 4910
rect 63870 4834 63922 4846
rect 66558 4898 66610 4910
rect 66558 4834 66610 4846
rect 69246 4898 69298 4910
rect 154814 4898 154866 4910
rect 136434 4846 136446 4898
rect 136498 4846 136510 4898
rect 140802 4846 140814 4898
rect 140866 4846 140878 4898
rect 146850 4846 146862 4898
rect 146914 4846 146926 4898
rect 69246 4834 69298 4846
rect 154814 4834 154866 4846
rect 155038 4898 155090 4910
rect 155038 4834 155090 4846
rect 156494 4898 156546 4910
rect 156494 4834 156546 4846
rect 158062 4898 158114 4910
rect 158062 4834 158114 4846
rect 160862 4898 160914 4910
rect 165342 4898 165394 4910
rect 164434 4846 164446 4898
rect 164498 4846 164510 4898
rect 160862 4834 160914 4846
rect 165342 4834 165394 4846
rect 165454 4898 165506 4910
rect 165454 4834 165506 4846
rect 166350 4898 166402 4910
rect 166350 4834 166402 4846
rect 166910 4898 166962 4910
rect 166910 4834 166962 4846
rect 1344 4730 218624 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 50558 4730
rect 50610 4678 50662 4730
rect 50714 4678 50766 4730
rect 50818 4678 81278 4730
rect 81330 4678 81382 4730
rect 81434 4678 81486 4730
rect 81538 4678 111998 4730
rect 112050 4678 112102 4730
rect 112154 4678 112206 4730
rect 112258 4678 142718 4730
rect 142770 4678 142822 4730
rect 142874 4678 142926 4730
rect 142978 4678 173438 4730
rect 173490 4678 173542 4730
rect 173594 4678 173646 4730
rect 173698 4678 204158 4730
rect 204210 4678 204262 4730
rect 204314 4678 204366 4730
rect 204418 4678 218624 4730
rect 1344 4644 218624 4678
rect 33182 4562 33234 4574
rect 33182 4498 33234 4510
rect 35646 4562 35698 4574
rect 35646 4498 35698 4510
rect 44494 4562 44546 4574
rect 44494 4498 44546 4510
rect 46958 4562 47010 4574
rect 46958 4498 47010 4510
rect 88062 4562 88114 4574
rect 88062 4498 88114 4510
rect 88958 4562 89010 4574
rect 149662 4562 149714 4574
rect 139234 4510 139246 4562
rect 139298 4510 139310 4562
rect 145170 4510 145182 4562
rect 145234 4510 145246 4562
rect 149090 4510 149102 4562
rect 149154 4510 149166 4562
rect 88958 4498 89010 4510
rect 149662 4498 149714 4510
rect 149886 4562 149938 4574
rect 151006 4562 151058 4574
rect 150658 4510 150670 4562
rect 150722 4510 150734 4562
rect 149886 4498 149938 4510
rect 151006 4498 151058 4510
rect 155038 4562 155090 4574
rect 155038 4498 155090 4510
rect 155262 4562 155314 4574
rect 155262 4498 155314 4510
rect 155374 4562 155426 4574
rect 155374 4498 155426 4510
rect 160862 4562 160914 4574
rect 160862 4498 160914 4510
rect 161422 4562 161474 4574
rect 161422 4498 161474 4510
rect 163662 4562 163714 4574
rect 163662 4498 163714 4510
rect 163774 4562 163826 4574
rect 163774 4498 163826 4510
rect 52558 4450 52610 4462
rect 150110 4450 150162 4462
rect 138786 4398 138798 4450
rect 138850 4398 138862 4450
rect 144946 4398 144958 4450
rect 145010 4398 145022 4450
rect 52558 4386 52610 4398
rect 150110 4386 150162 4398
rect 150222 4450 150274 4462
rect 155822 4450 155874 4462
rect 162766 4450 162818 4462
rect 152786 4398 152798 4450
rect 152850 4398 152862 4450
rect 153682 4398 153694 4450
rect 153746 4398 153758 4450
rect 156482 4398 156494 4450
rect 156546 4398 156558 4450
rect 150222 4386 150274 4398
rect 155822 4386 155874 4398
rect 162766 4386 162818 4398
rect 164222 4450 164274 4462
rect 164222 4386 164274 4398
rect 79550 4338 79602 4350
rect 5954 4286 5966 4338
rect 6018 4286 6030 4338
rect 32498 4286 32510 4338
rect 32562 4286 32574 4338
rect 44034 4286 44046 4338
rect 44098 4286 44110 4338
rect 51986 4286 51998 4338
rect 52050 4286 52062 4338
rect 57586 4286 57598 4338
rect 57650 4286 57662 4338
rect 68338 4286 68350 4338
rect 68402 4286 68414 4338
rect 78866 4286 78878 4338
rect 78930 4286 78942 4338
rect 79550 4274 79602 4286
rect 81342 4338 81394 4350
rect 149438 4338 149490 4350
rect 87042 4286 87054 4338
rect 87106 4286 87118 4338
rect 137330 4286 137342 4338
rect 137394 4286 137406 4338
rect 140242 4286 140254 4338
rect 140306 4286 140318 4338
rect 140466 4286 140478 4338
rect 140530 4286 140542 4338
rect 140914 4286 140926 4338
rect 140978 4286 140990 4338
rect 142258 4286 142270 4338
rect 142322 4286 142334 4338
rect 143490 4286 143502 4338
rect 143554 4286 143566 4338
rect 146066 4286 146078 4338
rect 146130 4286 146142 4338
rect 146626 4286 146638 4338
rect 146690 4286 146702 4338
rect 147074 4286 147086 4338
rect 147138 4286 147150 4338
rect 148418 4286 148430 4338
rect 148482 4286 148494 4338
rect 148866 4286 148878 4338
rect 148930 4286 148942 4338
rect 81342 4274 81394 4286
rect 149438 4274 149490 4286
rect 151454 4338 151506 4350
rect 161982 4338 162034 4350
rect 154578 4286 154590 4338
rect 154642 4286 154654 4338
rect 155586 4286 155598 4338
rect 155650 4286 155662 4338
rect 156258 4286 156270 4338
rect 156322 4286 156334 4338
rect 161634 4286 161646 4338
rect 161698 4286 161710 4338
rect 151454 4274 151506 4286
rect 161982 4274 162034 4286
rect 162206 4338 162258 4350
rect 162206 4274 162258 4286
rect 162430 4338 162482 4350
rect 162978 4286 162990 4338
rect 163042 4286 163054 4338
rect 163986 4286 163998 4338
rect 164050 4286 164062 4338
rect 162430 4274 162482 4286
rect 130846 4226 130898 4238
rect 130846 4162 130898 4174
rect 131294 4226 131346 4238
rect 131294 4162 131346 4174
rect 133758 4226 133810 4238
rect 133758 4162 133810 4174
rect 135326 4226 135378 4238
rect 135326 4162 135378 4174
rect 143054 4226 143106 4238
rect 165678 4226 165730 4238
rect 151218 4174 151230 4226
rect 151282 4174 151294 4226
rect 143054 4162 143106 4174
rect 165678 4162 165730 4174
rect 4062 4114 4114 4126
rect 41694 4114 41746 4126
rect 30594 4062 30606 4114
rect 30658 4062 30670 4114
rect 4062 4050 4114 4062
rect 41694 4050 41746 4062
rect 49758 4114 49810 4126
rect 49758 4050 49810 4062
rect 58606 4114 58658 4126
rect 58606 4050 58658 4062
rect 69358 4114 69410 4126
rect 69358 4050 69410 4062
rect 76638 4114 76690 4126
rect 76638 4050 76690 4062
rect 84702 4114 84754 4126
rect 84702 4050 84754 4062
rect 161758 4114 161810 4126
rect 163314 4062 163326 4114
rect 163378 4062 163390 4114
rect 161758 4050 161810 4062
rect 1344 3946 218624 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 65918 3946
rect 65970 3894 66022 3946
rect 66074 3894 66126 3946
rect 66178 3894 96638 3946
rect 96690 3894 96742 3946
rect 96794 3894 96846 3946
rect 96898 3894 127358 3946
rect 127410 3894 127462 3946
rect 127514 3894 127566 3946
rect 127618 3894 158078 3946
rect 158130 3894 158182 3946
rect 158234 3894 158286 3946
rect 158338 3894 188798 3946
rect 188850 3894 188902 3946
rect 188954 3894 189006 3946
rect 189058 3894 218624 3946
rect 1344 3860 218624 3894
rect 147858 3726 147870 3778
rect 147922 3775 147934 3778
rect 148754 3775 148766 3778
rect 147922 3729 148766 3775
rect 147922 3726 147934 3729
rect 148754 3726 148766 3729
rect 148818 3726 148830 3778
rect 161522 3726 161534 3778
rect 161586 3775 161598 3778
rect 162306 3775 162318 3778
rect 161586 3729 162318 3775
rect 161586 3726 161598 3729
rect 162306 3726 162318 3729
rect 162370 3726 162382 3778
rect 28590 3666 28642 3678
rect 28590 3602 28642 3614
rect 31502 3666 31554 3678
rect 36318 3666 36370 3678
rect 33170 3614 33182 3666
rect 33234 3614 33246 3666
rect 31502 3602 31554 3614
rect 36318 3602 36370 3614
rect 39230 3666 39282 3678
rect 39230 3602 39282 3614
rect 42926 3666 42978 3678
rect 42926 3602 42978 3614
rect 44382 3666 44434 3678
rect 44382 3602 44434 3614
rect 47630 3666 47682 3678
rect 47630 3602 47682 3614
rect 50542 3666 50594 3678
rect 50542 3602 50594 3614
rect 52894 3666 52946 3678
rect 52894 3602 52946 3614
rect 56030 3666 56082 3678
rect 56030 3602 56082 3614
rect 60510 3666 60562 3678
rect 60510 3602 60562 3614
rect 63982 3666 64034 3678
rect 63982 3602 64034 3614
rect 67454 3666 67506 3678
rect 67454 3602 67506 3614
rect 74286 3666 74338 3678
rect 74286 3602 74338 3614
rect 77198 3666 77250 3678
rect 82014 3666 82066 3678
rect 78866 3614 78878 3666
rect 78930 3614 78942 3666
rect 77198 3602 77250 3614
rect 82014 3602 82066 3614
rect 142830 3666 142882 3678
rect 142830 3602 142882 3614
rect 147422 3666 147474 3678
rect 147422 3602 147474 3614
rect 147870 3666 147922 3678
rect 147870 3602 147922 3614
rect 148318 3666 148370 3678
rect 148318 3602 148370 3614
rect 150334 3666 150386 3678
rect 150334 3602 150386 3614
rect 152798 3666 152850 3678
rect 156158 3666 156210 3678
rect 154466 3614 154478 3666
rect 154530 3614 154542 3666
rect 152798 3602 152850 3614
rect 156158 3602 156210 3614
rect 162318 3666 162370 3678
rect 211586 3614 211598 3666
rect 211650 3614 211662 3666
rect 213938 3614 213950 3666
rect 214002 3614 214014 3666
rect 216626 3614 216638 3666
rect 216690 3614 216702 3666
rect 162318 3602 162370 3614
rect 148766 3554 148818 3566
rect 151342 3554 151394 3566
rect 30930 3502 30942 3554
rect 30994 3502 31006 3554
rect 35410 3502 35422 3554
rect 35474 3502 35486 3554
rect 38658 3502 38670 3554
rect 38722 3502 38734 3554
rect 42354 3502 42366 3554
rect 42418 3502 42430 3554
rect 46722 3502 46734 3554
rect 46786 3502 46798 3554
rect 49970 3502 49982 3554
rect 50034 3502 50046 3554
rect 51874 3502 51886 3554
rect 51938 3502 51950 3554
rect 55010 3502 55022 3554
rect 55074 3502 55086 3554
rect 59490 3502 59502 3554
rect 59554 3502 59566 3554
rect 62962 3502 62974 3554
rect 63026 3502 63038 3554
rect 66434 3502 66446 3554
rect 66498 3502 66510 3554
rect 70914 3502 70926 3554
rect 70978 3502 70990 3554
rect 76514 3502 76526 3554
rect 76578 3502 76590 3554
rect 81106 3502 81118 3554
rect 81170 3502 81182 3554
rect 84354 3502 84366 3554
rect 84418 3502 84430 3554
rect 88722 3502 88734 3554
rect 88786 3502 88798 3554
rect 150882 3502 150894 3554
rect 150946 3502 150958 3554
rect 148766 3490 148818 3502
rect 151342 3490 151394 3502
rect 152014 3554 152066 3566
rect 152014 3490 152066 3502
rect 152238 3554 152290 3566
rect 152238 3490 152290 3502
rect 152462 3554 152514 3566
rect 152462 3490 152514 3502
rect 152686 3554 152738 3566
rect 152686 3490 152738 3502
rect 153358 3554 153410 3566
rect 153358 3490 153410 3502
rect 154030 3554 154082 3566
rect 155710 3554 155762 3566
rect 155026 3502 155038 3554
rect 155090 3502 155102 3554
rect 154030 3490 154082 3502
rect 155710 3490 155762 3502
rect 162654 3554 162706 3566
rect 197934 3554 197986 3566
rect 165666 3502 165678 3554
rect 165730 3502 165742 3554
rect 170706 3502 170718 3554
rect 170770 3502 170782 3554
rect 176082 3502 176094 3554
rect 176146 3502 176158 3554
rect 178770 3502 178782 3554
rect 178834 3502 178846 3554
rect 184706 3502 184718 3554
rect 184770 3502 184782 3554
rect 186834 3502 186846 3554
rect 186898 3502 186910 3554
rect 189522 3502 189534 3554
rect 189586 3502 189598 3554
rect 192322 3502 192334 3554
rect 192386 3502 192398 3554
rect 162654 3490 162706 3502
rect 197934 3490 197986 3502
rect 205998 3554 206050 3566
rect 205998 3490 206050 3502
rect 84926 3442 84978 3454
rect 89630 3442 89682 3454
rect 40562 3390 40574 3442
rect 40626 3390 40638 3442
rect 86930 3390 86942 3442
rect 86994 3390 87006 3442
rect 84926 3378 84978 3390
rect 89630 3378 89682 3390
rect 89854 3442 89906 3454
rect 92654 3442 92706 3454
rect 90178 3390 90190 3442
rect 90242 3390 90254 3442
rect 89854 3378 89906 3390
rect 92654 3378 92706 3390
rect 93102 3442 93154 3454
rect 95006 3442 95058 3454
rect 93426 3390 93438 3442
rect 93490 3390 93502 3442
rect 93102 3378 93154 3390
rect 95006 3378 95058 3390
rect 95230 3442 95282 3454
rect 97694 3442 97746 3454
rect 95554 3390 95566 3442
rect 95618 3390 95630 3442
rect 95230 3378 95282 3390
rect 97694 3378 97746 3390
rect 97918 3442 97970 3454
rect 97918 3378 97970 3390
rect 98254 3442 98306 3454
rect 98254 3378 98306 3390
rect 100270 3442 100322 3454
rect 100270 3378 100322 3390
rect 100718 3442 100770 3454
rect 100718 3378 100770 3390
rect 101054 3442 101106 3454
rect 101054 3378 101106 3390
rect 103070 3442 103122 3454
rect 103070 3378 103122 3390
rect 103294 3442 103346 3454
rect 103294 3378 103346 3390
rect 103630 3442 103682 3454
rect 103630 3378 103682 3390
rect 105758 3442 105810 3454
rect 105758 3378 105810 3390
rect 105982 3442 106034 3454
rect 105982 3378 106034 3390
rect 106318 3442 106370 3454
rect 106318 3378 106370 3390
rect 107886 3442 107938 3454
rect 107886 3378 107938 3390
rect 108670 3442 108722 3454
rect 108670 3378 108722 3390
rect 109006 3442 109058 3454
rect 109006 3378 109058 3390
rect 111694 3442 111746 3454
rect 111694 3378 111746 3390
rect 112142 3442 112194 3454
rect 113822 3442 113874 3454
rect 112466 3390 112478 3442
rect 112530 3390 112542 3442
rect 112142 3378 112194 3390
rect 113822 3378 113874 3390
rect 114046 3442 114098 3454
rect 114046 3378 114098 3390
rect 114382 3442 114434 3454
rect 114382 3378 114434 3390
rect 116510 3442 116562 3454
rect 116510 3378 116562 3390
rect 116734 3442 116786 3454
rect 116734 3378 116786 3390
rect 117070 3442 117122 3454
rect 117070 3378 117122 3390
rect 119310 3442 119362 3454
rect 119310 3378 119362 3390
rect 119758 3442 119810 3454
rect 119758 3378 119810 3390
rect 120094 3442 120146 3454
rect 120094 3378 120146 3390
rect 121886 3442 121938 3454
rect 121886 3378 121938 3390
rect 122110 3442 122162 3454
rect 122110 3378 122162 3390
rect 124574 3442 124626 3454
rect 124574 3378 124626 3390
rect 124798 3442 124850 3454
rect 126926 3442 126978 3454
rect 125122 3390 125134 3442
rect 125186 3390 125198 3442
rect 124798 3378 124850 3390
rect 126926 3378 126978 3390
rect 127486 3442 127538 3454
rect 127486 3378 127538 3390
rect 127822 3442 127874 3454
rect 127822 3378 127874 3390
rect 129950 3442 130002 3454
rect 129950 3378 130002 3390
rect 130174 3442 130226 3454
rect 130174 3378 130226 3390
rect 130510 3442 130562 3454
rect 130510 3378 130562 3390
rect 132638 3442 132690 3454
rect 132638 3378 132690 3390
rect 132862 3442 132914 3454
rect 135326 3442 135378 3454
rect 133186 3390 133198 3442
rect 133250 3390 133262 3442
rect 132862 3378 132914 3390
rect 135326 3378 135378 3390
rect 135550 3442 135602 3454
rect 138350 3442 138402 3454
rect 135874 3390 135886 3442
rect 135938 3390 135950 3442
rect 135550 3378 135602 3390
rect 138350 3378 138402 3390
rect 138798 3442 138850 3454
rect 140702 3442 140754 3454
rect 139122 3390 139134 3442
rect 139186 3390 139198 3442
rect 138798 3378 138850 3390
rect 140702 3378 140754 3390
rect 140926 3442 140978 3454
rect 140926 3378 140978 3390
rect 141262 3442 141314 3454
rect 141262 3378 141314 3390
rect 143390 3442 143442 3454
rect 143390 3378 143442 3390
rect 143614 3442 143666 3454
rect 143614 3378 143666 3390
rect 143950 3442 144002 3454
rect 143950 3378 144002 3390
rect 145966 3442 146018 3454
rect 145966 3378 146018 3390
rect 146414 3442 146466 3454
rect 146414 3378 146466 3390
rect 146750 3442 146802 3454
rect 146750 3378 146802 3390
rect 148990 3442 149042 3454
rect 155262 3442 155314 3454
rect 149314 3390 149326 3442
rect 149378 3390 149390 3442
rect 153010 3390 153022 3442
rect 153074 3390 153086 3442
rect 148990 3378 149042 3390
rect 155262 3378 155314 3390
rect 156606 3442 156658 3454
rect 156606 3378 156658 3390
rect 157390 3442 157442 3454
rect 157390 3378 157442 3390
rect 157838 3442 157890 3454
rect 157838 3378 157890 3390
rect 158174 3442 158226 3454
rect 158174 3378 158226 3390
rect 159518 3442 159570 3454
rect 159518 3378 159570 3390
rect 160078 3442 160130 3454
rect 160078 3378 160130 3390
rect 161982 3442 162034 3454
rect 163326 3442 163378 3454
rect 162978 3390 162990 3442
rect 163042 3390 163054 3442
rect 161982 3378 162034 3390
rect 163326 3378 163378 3390
rect 163662 3442 163714 3454
rect 163662 3378 163714 3390
rect 165006 3442 165058 3454
rect 165006 3378 165058 3390
rect 165454 3442 165506 3454
rect 165454 3378 165506 3390
rect 167582 3442 167634 3454
rect 167582 3378 167634 3390
rect 168142 3442 168194 3454
rect 168142 3378 168194 3390
rect 170270 3442 170322 3454
rect 170270 3378 170322 3390
rect 172622 3442 172674 3454
rect 172622 3378 172674 3390
rect 173182 3442 173234 3454
rect 173182 3378 173234 3390
rect 173518 3442 173570 3454
rect 173518 3378 173570 3390
rect 175646 3442 175698 3454
rect 175646 3378 175698 3390
rect 178334 3442 178386 3454
rect 178334 3378 178386 3390
rect 181022 3442 181074 3454
rect 181022 3378 181074 3390
rect 181582 3442 181634 3454
rect 181582 3378 181634 3390
rect 184046 3442 184098 3454
rect 184046 3378 184098 3390
rect 186398 3442 186450 3454
rect 186398 3378 186450 3390
rect 189086 3442 189138 3454
rect 189086 3378 189138 3390
rect 191662 3442 191714 3454
rect 191662 3378 191714 3390
rect 194462 3442 194514 3454
rect 194462 3378 194514 3390
rect 195022 3442 195074 3454
rect 195022 3378 195074 3390
rect 197150 3442 197202 3454
rect 197150 3378 197202 3390
rect 197374 3442 197426 3454
rect 197374 3378 197426 3390
rect 199278 3442 199330 3454
rect 199278 3378 199330 3390
rect 200062 3442 200114 3454
rect 200062 3378 200114 3390
rect 200622 3442 200674 3454
rect 200622 3378 200674 3390
rect 203086 3442 203138 3454
rect 203086 3378 203138 3390
rect 203534 3442 203586 3454
rect 203534 3378 203586 3390
rect 204094 3442 204146 3454
rect 204094 3378 204146 3390
rect 205214 3442 205266 3454
rect 205214 3378 205266 3390
rect 205438 3442 205490 3454
rect 205438 3378 205490 3390
rect 207902 3442 207954 3454
rect 207902 3378 207954 3390
rect 208126 3442 208178 3454
rect 208126 3378 208178 3390
rect 208686 3442 208738 3454
rect 208686 3378 208738 3390
rect 210702 3442 210754 3454
rect 210702 3378 210754 3390
rect 211150 3442 211202 3454
rect 211150 3378 211202 3390
rect 213278 3442 213330 3454
rect 213278 3378 213330 3390
rect 213502 3442 213554 3454
rect 213502 3378 213554 3390
rect 215966 3442 216018 3454
rect 215966 3378 216018 3390
rect 216190 3442 216242 3454
rect 216190 3378 216242 3390
rect 6526 3330 6578 3342
rect 6526 3266 6578 3278
rect 9326 3330 9378 3342
rect 9326 3266 9378 3278
rect 11902 3330 11954 3342
rect 11902 3266 11954 3278
rect 14590 3330 14642 3342
rect 14590 3266 14642 3278
rect 17278 3330 17330 3342
rect 17278 3266 17330 3278
rect 19966 3330 20018 3342
rect 19966 3266 20018 3278
rect 22654 3330 22706 3342
rect 22654 3266 22706 3278
rect 25342 3330 25394 3342
rect 25342 3266 25394 3278
rect 71934 3330 71986 3342
rect 71934 3266 71986 3278
rect 122446 3330 122498 3342
rect 122446 3266 122498 3278
rect 159742 3330 159794 3342
rect 159742 3266 159794 3278
rect 167806 3330 167858 3342
rect 167806 3266 167858 3278
rect 170494 3330 170546 3342
rect 170494 3266 170546 3278
rect 175870 3330 175922 3342
rect 175870 3266 175922 3278
rect 178558 3330 178610 3342
rect 178558 3266 178610 3278
rect 181246 3330 181298 3342
rect 181246 3266 181298 3278
rect 184494 3330 184546 3342
rect 184494 3266 184546 3278
rect 186622 3330 186674 3342
rect 186622 3266 186674 3278
rect 189310 3330 189362 3342
rect 189310 3266 189362 3278
rect 192110 3330 192162 3342
rect 192110 3266 192162 3278
rect 194686 3330 194738 3342
rect 194686 3266 194738 3278
rect 1344 3162 218624 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 50558 3162
rect 50610 3110 50662 3162
rect 50714 3110 50766 3162
rect 50818 3110 81278 3162
rect 81330 3110 81382 3162
rect 81434 3110 81486 3162
rect 81538 3110 111998 3162
rect 112050 3110 112102 3162
rect 112154 3110 112206 3162
rect 112258 3110 142718 3162
rect 142770 3110 142822 3162
rect 142874 3110 142926 3162
rect 142978 3110 173438 3162
rect 173490 3110 173542 3162
rect 173594 3110 173646 3162
rect 173698 3110 204158 3162
rect 204210 3110 204262 3162
rect 204314 3110 204366 3162
rect 204418 3110 218624 3162
rect 1344 3076 218624 3110
<< via1 >>
rect 27134 46398 27186 46450
rect 27806 46398 27858 46450
rect 28366 46398 28418 46450
rect 168702 46398 168754 46450
rect 169486 46398 169538 46450
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 65918 46230 65970 46282
rect 66022 46230 66074 46282
rect 66126 46230 66178 46282
rect 96638 46230 96690 46282
rect 96742 46230 96794 46282
rect 96846 46230 96898 46282
rect 127358 46230 127410 46282
rect 127462 46230 127514 46282
rect 127566 46230 127618 46282
rect 158078 46230 158130 46282
rect 158182 46230 158234 46282
rect 158286 46230 158338 46282
rect 188798 46230 188850 46282
rect 188902 46230 188954 46282
rect 189006 46230 189058 46282
rect 47742 46062 47794 46114
rect 51774 46062 51826 46114
rect 55806 46062 55858 46114
rect 59726 46062 59778 46114
rect 63534 46062 63586 46114
rect 150446 46062 150498 46114
rect 6974 45950 7026 46002
rect 11006 45950 11058 46002
rect 15038 45950 15090 46002
rect 19070 45950 19122 46002
rect 23102 45950 23154 46002
rect 27806 45950 27858 46002
rect 31614 45950 31666 46002
rect 35422 45950 35474 46002
rect 39230 45950 39282 46002
rect 40238 45950 40290 46002
rect 43150 45950 43202 46002
rect 67454 45950 67506 46002
rect 71486 45950 71538 46002
rect 79550 45950 79602 46002
rect 83582 45950 83634 46002
rect 87614 45950 87666 46002
rect 91646 45950 91698 46002
rect 95678 45950 95730 46002
rect 100158 45950 100210 46002
rect 103966 45950 104018 46002
rect 107774 45950 107826 46002
rect 111694 45950 111746 46002
rect 115502 45950 115554 46002
rect 119310 45950 119362 46002
rect 123902 45950 123954 46002
rect 127934 45950 127986 46002
rect 131966 45950 132018 46002
rect 135998 45950 136050 46002
rect 140030 45950 140082 46002
rect 144062 45950 144114 46002
rect 156158 45950 156210 46002
rect 160190 45950 160242 46002
rect 164222 45950 164274 46002
rect 168702 45950 168754 46002
rect 172510 45950 172562 46002
rect 176318 45950 176370 46002
rect 180238 45950 180290 46002
rect 184046 45950 184098 46002
rect 187854 45950 187906 46002
rect 192446 45950 192498 46002
rect 193118 45950 193170 46002
rect 196478 45950 196530 46002
rect 200510 45950 200562 46002
rect 204542 45950 204594 46002
rect 205214 45950 205266 46002
rect 208574 45950 208626 46002
rect 212606 45950 212658 46002
rect 216638 45950 216690 46002
rect 217534 45950 217586 46002
rect 7422 45838 7474 45890
rect 11230 45838 11282 45890
rect 15262 45838 15314 45890
rect 15822 45838 15874 45890
rect 19294 45838 19346 45890
rect 19854 45838 19906 45890
rect 23326 45838 23378 45890
rect 23886 45838 23938 45890
rect 28366 45838 28418 45890
rect 28926 45838 28978 45890
rect 32174 45838 32226 45890
rect 32734 45838 32786 45890
rect 35982 45838 36034 45890
rect 36542 45838 36594 45890
rect 39790 45838 39842 45890
rect 43598 45838 43650 45890
rect 44158 45838 44210 45890
rect 50094 45838 50146 45890
rect 54126 45838 54178 45890
rect 55134 45838 55186 45890
rect 58158 45838 58210 45890
rect 62078 45838 62130 45890
rect 65886 45838 65938 45890
rect 69694 45838 69746 45890
rect 73502 45838 73554 45890
rect 79774 45838 79826 45890
rect 83806 45838 83858 45890
rect 87838 45838 87890 45890
rect 91870 45838 91922 45890
rect 95902 45838 95954 45890
rect 100830 45838 100882 45890
rect 104638 45838 104690 45890
rect 108334 45838 108386 45890
rect 112142 45838 112194 45890
rect 116062 45838 116114 45890
rect 120094 45838 120146 45890
rect 124126 45838 124178 45890
rect 128158 45838 128210 45890
rect 132190 45838 132242 45890
rect 136446 45838 136498 45890
rect 140478 45838 140530 45890
rect 144510 45838 144562 45890
rect 152798 45838 152850 45890
rect 156382 45838 156434 45890
rect 160638 45838 160690 45890
rect 164670 45838 164722 45890
rect 169486 45838 169538 45890
rect 173294 45838 173346 45890
rect 177102 45838 177154 45890
rect 180910 45838 180962 45890
rect 184830 45838 184882 45890
rect 188638 45838 188690 45890
rect 192670 45838 192722 45890
rect 196702 45838 196754 45890
rect 200734 45838 200786 45890
rect 204766 45838 204818 45890
rect 208798 45838 208850 45890
rect 212830 45838 212882 45890
rect 216862 45838 216914 45890
rect 12350 45726 12402 45778
rect 66558 45726 66610 45778
rect 189198 45726 189250 45778
rect 197262 45726 197314 45778
rect 201294 45726 201346 45778
rect 209358 45726 209410 45778
rect 213950 45726 214002 45778
rect 7198 45614 7250 45666
rect 50542 45614 50594 45666
rect 58942 45614 58994 45666
rect 62750 45614 62802 45666
rect 70366 45614 70418 45666
rect 74174 45614 74226 45666
rect 80110 45614 80162 45666
rect 84142 45614 84194 45666
rect 88174 45614 88226 45666
rect 92206 45614 92258 45666
rect 96238 45614 96290 45666
rect 101054 45614 101106 45666
rect 104862 45614 104914 45666
rect 108670 45614 108722 45666
rect 112478 45614 112530 45666
rect 116398 45614 116450 45666
rect 120430 45614 120482 45666
rect 124462 45614 124514 45666
rect 128494 45614 128546 45666
rect 132526 45614 132578 45666
rect 136222 45614 136274 45666
rect 140254 45614 140306 45666
rect 144286 45614 144338 45666
rect 153246 45614 153298 45666
rect 156718 45614 156770 45666
rect 160414 45614 160466 45666
rect 164446 45614 164498 45666
rect 169262 45614 169314 45666
rect 173070 45614 173122 45666
rect 176878 45614 176930 45666
rect 180686 45614 180738 45666
rect 184606 45614 184658 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 50558 45446 50610 45498
rect 50662 45446 50714 45498
rect 50766 45446 50818 45498
rect 81278 45446 81330 45498
rect 81382 45446 81434 45498
rect 81486 45446 81538 45498
rect 111998 45446 112050 45498
rect 112102 45446 112154 45498
rect 112206 45446 112258 45498
rect 142718 45446 142770 45498
rect 142822 45446 142874 45498
rect 142926 45446 142978 45498
rect 173438 45446 173490 45498
rect 173542 45446 173594 45498
rect 173646 45446 173698 45498
rect 204158 45446 204210 45498
rect 204262 45446 204314 45498
rect 204366 45446 204418 45498
rect 153358 45278 153410 45330
rect 140590 45166 140642 45218
rect 78318 45054 78370 45106
rect 78878 45054 78930 45106
rect 141598 45054 141650 45106
rect 152350 45054 152402 45106
rect 75966 44942 76018 44994
rect 135214 44942 135266 44994
rect 138126 44942 138178 44994
rect 138686 44942 138738 44994
rect 139694 44942 139746 44994
rect 139806 44942 139858 44994
rect 152126 44942 152178 44994
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 65918 44662 65970 44714
rect 66022 44662 66074 44714
rect 66126 44662 66178 44714
rect 96638 44662 96690 44714
rect 96742 44662 96794 44714
rect 96846 44662 96898 44714
rect 127358 44662 127410 44714
rect 127462 44662 127514 44714
rect 127566 44662 127618 44714
rect 158078 44662 158130 44714
rect 158182 44662 158234 44714
rect 158286 44662 158338 44714
rect 188798 44662 188850 44714
rect 188902 44662 188954 44714
rect 189006 44662 189058 44714
rect 132638 44382 132690 44434
rect 134766 44382 134818 44434
rect 135886 44382 135938 44434
rect 138014 44382 138066 44434
rect 139694 44382 139746 44434
rect 141822 44382 141874 44434
rect 131966 44270 132018 44322
rect 135102 44270 135154 44322
rect 138910 44270 138962 44322
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 50558 43878 50610 43930
rect 50662 43878 50714 43930
rect 50766 43878 50818 43930
rect 81278 43878 81330 43930
rect 81382 43878 81434 43930
rect 81486 43878 81538 43930
rect 111998 43878 112050 43930
rect 112102 43878 112154 43930
rect 112206 43878 112258 43930
rect 142718 43878 142770 43930
rect 142822 43878 142874 43930
rect 142926 43878 142978 43930
rect 173438 43878 173490 43930
rect 173542 43878 173594 43930
rect 173646 43878 173698 43930
rect 204158 43878 204210 43930
rect 204262 43878 204314 43930
rect 204366 43878 204418 43930
rect 135886 43598 135938 43650
rect 136110 43598 136162 43650
rect 139694 43598 139746 43650
rect 135774 43486 135826 43538
rect 136222 43486 136274 43538
rect 140366 43486 140418 43538
rect 135102 43374 135154 43426
rect 137230 43374 137282 43426
rect 137566 43374 137618 43426
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 65918 43094 65970 43146
rect 66022 43094 66074 43146
rect 66126 43094 66178 43146
rect 96638 43094 96690 43146
rect 96742 43094 96794 43146
rect 96846 43094 96898 43146
rect 127358 43094 127410 43146
rect 127462 43094 127514 43146
rect 127566 43094 127618 43146
rect 158078 43094 158130 43146
rect 158182 43094 158234 43146
rect 158286 43094 158338 43146
rect 188798 43094 188850 43146
rect 188902 43094 188954 43146
rect 189006 43094 189058 43146
rect 137790 42926 137842 42978
rect 138126 42926 138178 42978
rect 137902 42702 137954 42754
rect 137790 42478 137842 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 50558 42310 50610 42362
rect 50662 42310 50714 42362
rect 50766 42310 50818 42362
rect 81278 42310 81330 42362
rect 81382 42310 81434 42362
rect 81486 42310 81538 42362
rect 111998 42310 112050 42362
rect 112102 42310 112154 42362
rect 112206 42310 112258 42362
rect 142718 42310 142770 42362
rect 142822 42310 142874 42362
rect 142926 42310 142978 42362
rect 173438 42310 173490 42362
rect 173542 42310 173594 42362
rect 173646 42310 173698 42362
rect 204158 42310 204210 42362
rect 204262 42310 204314 42362
rect 204366 42310 204418 42362
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 65918 41526 65970 41578
rect 66022 41526 66074 41578
rect 66126 41526 66178 41578
rect 96638 41526 96690 41578
rect 96742 41526 96794 41578
rect 96846 41526 96898 41578
rect 127358 41526 127410 41578
rect 127462 41526 127514 41578
rect 127566 41526 127618 41578
rect 158078 41526 158130 41578
rect 158182 41526 158234 41578
rect 158286 41526 158338 41578
rect 188798 41526 188850 41578
rect 188902 41526 188954 41578
rect 189006 41526 189058 41578
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 50558 40742 50610 40794
rect 50662 40742 50714 40794
rect 50766 40742 50818 40794
rect 81278 40742 81330 40794
rect 81382 40742 81434 40794
rect 81486 40742 81538 40794
rect 111998 40742 112050 40794
rect 112102 40742 112154 40794
rect 112206 40742 112258 40794
rect 142718 40742 142770 40794
rect 142822 40742 142874 40794
rect 142926 40742 142978 40794
rect 173438 40742 173490 40794
rect 173542 40742 173594 40794
rect 173646 40742 173698 40794
rect 204158 40742 204210 40794
rect 204262 40742 204314 40794
rect 204366 40742 204418 40794
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 65918 39958 65970 40010
rect 66022 39958 66074 40010
rect 66126 39958 66178 40010
rect 96638 39958 96690 40010
rect 96742 39958 96794 40010
rect 96846 39958 96898 40010
rect 127358 39958 127410 40010
rect 127462 39958 127514 40010
rect 127566 39958 127618 40010
rect 158078 39958 158130 40010
rect 158182 39958 158234 40010
rect 158286 39958 158338 40010
rect 188798 39958 188850 40010
rect 188902 39958 188954 40010
rect 189006 39958 189058 40010
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 50558 39174 50610 39226
rect 50662 39174 50714 39226
rect 50766 39174 50818 39226
rect 81278 39174 81330 39226
rect 81382 39174 81434 39226
rect 81486 39174 81538 39226
rect 111998 39174 112050 39226
rect 112102 39174 112154 39226
rect 112206 39174 112258 39226
rect 142718 39174 142770 39226
rect 142822 39174 142874 39226
rect 142926 39174 142978 39226
rect 173438 39174 173490 39226
rect 173542 39174 173594 39226
rect 173646 39174 173698 39226
rect 204158 39174 204210 39226
rect 204262 39174 204314 39226
rect 204366 39174 204418 39226
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 65918 38390 65970 38442
rect 66022 38390 66074 38442
rect 66126 38390 66178 38442
rect 96638 38390 96690 38442
rect 96742 38390 96794 38442
rect 96846 38390 96898 38442
rect 127358 38390 127410 38442
rect 127462 38390 127514 38442
rect 127566 38390 127618 38442
rect 158078 38390 158130 38442
rect 158182 38390 158234 38442
rect 158286 38390 158338 38442
rect 188798 38390 188850 38442
rect 188902 38390 188954 38442
rect 189006 38390 189058 38442
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 50558 37606 50610 37658
rect 50662 37606 50714 37658
rect 50766 37606 50818 37658
rect 81278 37606 81330 37658
rect 81382 37606 81434 37658
rect 81486 37606 81538 37658
rect 111998 37606 112050 37658
rect 112102 37606 112154 37658
rect 112206 37606 112258 37658
rect 142718 37606 142770 37658
rect 142822 37606 142874 37658
rect 142926 37606 142978 37658
rect 173438 37606 173490 37658
rect 173542 37606 173594 37658
rect 173646 37606 173698 37658
rect 204158 37606 204210 37658
rect 204262 37606 204314 37658
rect 204366 37606 204418 37658
rect 119310 37214 119362 37266
rect 118750 37102 118802 37154
rect 124238 37102 124290 37154
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 65918 36822 65970 36874
rect 66022 36822 66074 36874
rect 66126 36822 66178 36874
rect 96638 36822 96690 36874
rect 96742 36822 96794 36874
rect 96846 36822 96898 36874
rect 127358 36822 127410 36874
rect 127462 36822 127514 36874
rect 127566 36822 127618 36874
rect 158078 36822 158130 36874
rect 158182 36822 158234 36874
rect 158286 36822 158338 36874
rect 188798 36822 188850 36874
rect 188902 36822 188954 36874
rect 189006 36822 189058 36874
rect 131070 36430 131122 36482
rect 135998 36318 136050 36370
rect 130510 36206 130562 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 50558 36038 50610 36090
rect 50662 36038 50714 36090
rect 50766 36038 50818 36090
rect 81278 36038 81330 36090
rect 81382 36038 81434 36090
rect 81486 36038 81538 36090
rect 111998 36038 112050 36090
rect 112102 36038 112154 36090
rect 112206 36038 112258 36090
rect 142718 36038 142770 36090
rect 142822 36038 142874 36090
rect 142926 36038 142978 36090
rect 173438 36038 173490 36090
rect 173542 36038 173594 36090
rect 173646 36038 173698 36090
rect 204158 36038 204210 36090
rect 204262 36038 204314 36090
rect 204366 36038 204418 36090
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 65918 35254 65970 35306
rect 66022 35254 66074 35306
rect 66126 35254 66178 35306
rect 96638 35254 96690 35306
rect 96742 35254 96794 35306
rect 96846 35254 96898 35306
rect 127358 35254 127410 35306
rect 127462 35254 127514 35306
rect 127566 35254 127618 35306
rect 158078 35254 158130 35306
rect 158182 35254 158234 35306
rect 158286 35254 158338 35306
rect 188798 35254 188850 35306
rect 188902 35254 188954 35306
rect 189006 35254 189058 35306
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 50558 34470 50610 34522
rect 50662 34470 50714 34522
rect 50766 34470 50818 34522
rect 81278 34470 81330 34522
rect 81382 34470 81434 34522
rect 81486 34470 81538 34522
rect 111998 34470 112050 34522
rect 112102 34470 112154 34522
rect 112206 34470 112258 34522
rect 142718 34470 142770 34522
rect 142822 34470 142874 34522
rect 142926 34470 142978 34522
rect 173438 34470 173490 34522
rect 173542 34470 173594 34522
rect 173646 34470 173698 34522
rect 204158 34470 204210 34522
rect 204262 34470 204314 34522
rect 204366 34470 204418 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 65918 33686 65970 33738
rect 66022 33686 66074 33738
rect 66126 33686 66178 33738
rect 96638 33686 96690 33738
rect 96742 33686 96794 33738
rect 96846 33686 96898 33738
rect 127358 33686 127410 33738
rect 127462 33686 127514 33738
rect 127566 33686 127618 33738
rect 158078 33686 158130 33738
rect 158182 33686 158234 33738
rect 158286 33686 158338 33738
rect 188798 33686 188850 33738
rect 188902 33686 188954 33738
rect 189006 33686 189058 33738
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 50558 32902 50610 32954
rect 50662 32902 50714 32954
rect 50766 32902 50818 32954
rect 81278 32902 81330 32954
rect 81382 32902 81434 32954
rect 81486 32902 81538 32954
rect 111998 32902 112050 32954
rect 112102 32902 112154 32954
rect 112206 32902 112258 32954
rect 142718 32902 142770 32954
rect 142822 32902 142874 32954
rect 142926 32902 142978 32954
rect 173438 32902 173490 32954
rect 173542 32902 173594 32954
rect 173646 32902 173698 32954
rect 204158 32902 204210 32954
rect 204262 32902 204314 32954
rect 204366 32902 204418 32954
rect 117182 32734 117234 32786
rect 116734 32510 116786 32562
rect 112590 32398 112642 32450
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 65918 32118 65970 32170
rect 66022 32118 66074 32170
rect 66126 32118 66178 32170
rect 96638 32118 96690 32170
rect 96742 32118 96794 32170
rect 96846 32118 96898 32170
rect 127358 32118 127410 32170
rect 127462 32118 127514 32170
rect 127566 32118 127618 32170
rect 158078 32118 158130 32170
rect 158182 32118 158234 32170
rect 158286 32118 158338 32170
rect 188798 32118 188850 32170
rect 188902 32118 188954 32170
rect 189006 32118 189058 32170
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 50558 31334 50610 31386
rect 50662 31334 50714 31386
rect 50766 31334 50818 31386
rect 81278 31334 81330 31386
rect 81382 31334 81434 31386
rect 81486 31334 81538 31386
rect 111998 31334 112050 31386
rect 112102 31334 112154 31386
rect 112206 31334 112258 31386
rect 142718 31334 142770 31386
rect 142822 31334 142874 31386
rect 142926 31334 142978 31386
rect 173438 31334 173490 31386
rect 173542 31334 173594 31386
rect 173646 31334 173698 31386
rect 204158 31334 204210 31386
rect 204262 31334 204314 31386
rect 204366 31334 204418 31386
rect 117294 31166 117346 31218
rect 108894 30942 108946 30994
rect 116734 30942 116786 30994
rect 137342 30942 137394 30994
rect 108222 30830 108274 30882
rect 109454 30830 109506 30882
rect 109902 30830 109954 30882
rect 113598 30830 113650 30882
rect 116062 30830 116114 30882
rect 136334 30830 136386 30882
rect 136782 30830 136834 30882
rect 138126 30830 138178 30882
rect 140254 30830 140306 30882
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 65918 30550 65970 30602
rect 66022 30550 66074 30602
rect 66126 30550 66178 30602
rect 96638 30550 96690 30602
rect 96742 30550 96794 30602
rect 96846 30550 96898 30602
rect 127358 30550 127410 30602
rect 127462 30550 127514 30602
rect 127566 30550 127618 30602
rect 158078 30550 158130 30602
rect 158182 30550 158234 30602
rect 158286 30550 158338 30602
rect 188798 30550 188850 30602
rect 188902 30550 188954 30602
rect 189006 30550 189058 30602
rect 113374 30270 113426 30322
rect 135774 30270 135826 30322
rect 96238 30158 96290 30210
rect 96686 30158 96738 30210
rect 104414 30158 104466 30210
rect 104974 30158 105026 30210
rect 112366 30158 112418 30210
rect 117630 30158 117682 30210
rect 117966 30158 118018 30210
rect 128942 30158 128994 30210
rect 129950 30158 130002 30210
rect 132638 30158 132690 30210
rect 132862 30158 132914 30210
rect 136222 30158 136274 30210
rect 95454 30046 95506 30098
rect 97134 30046 97186 30098
rect 103742 30046 103794 30098
rect 105422 30046 105474 30098
rect 111694 30046 111746 30098
rect 112926 30046 112978 30098
rect 118750 30046 118802 30098
rect 128270 30046 128322 30098
rect 129502 30046 129554 30098
rect 133646 30046 133698 30098
rect 121326 29934 121378 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 50558 29766 50610 29818
rect 50662 29766 50714 29818
rect 50766 29766 50818 29818
rect 81278 29766 81330 29818
rect 81382 29766 81434 29818
rect 81486 29766 81538 29818
rect 111998 29766 112050 29818
rect 112102 29766 112154 29818
rect 112206 29766 112258 29818
rect 142718 29766 142770 29818
rect 142822 29766 142874 29818
rect 142926 29766 142978 29818
rect 173438 29766 173490 29818
rect 173542 29766 173594 29818
rect 173646 29766 173698 29818
rect 204158 29766 204210 29818
rect 204262 29766 204314 29818
rect 204366 29766 204418 29818
rect 101278 29598 101330 29650
rect 125358 29598 125410 29650
rect 133982 29598 134034 29650
rect 134430 29598 134482 29650
rect 135774 29486 135826 29538
rect 100830 29374 100882 29426
rect 124462 29374 124514 29426
rect 134990 29374 135042 29426
rect 100046 29262 100098 29314
rect 101726 29262 101778 29314
rect 123678 29262 123730 29314
rect 124910 29262 124962 29314
rect 137902 29262 137954 29314
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 65918 28982 65970 29034
rect 66022 28982 66074 29034
rect 66126 28982 66178 29034
rect 96638 28982 96690 29034
rect 96742 28982 96794 29034
rect 96846 28982 96898 29034
rect 127358 28982 127410 29034
rect 127462 28982 127514 29034
rect 127566 28982 127618 29034
rect 158078 28982 158130 29034
rect 158182 28982 158234 29034
rect 158286 28982 158338 29034
rect 188798 28982 188850 29034
rect 188902 28982 188954 29034
rect 189006 28982 189058 29034
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 50558 28198 50610 28250
rect 50662 28198 50714 28250
rect 50766 28198 50818 28250
rect 81278 28198 81330 28250
rect 81382 28198 81434 28250
rect 81486 28198 81538 28250
rect 111998 28198 112050 28250
rect 112102 28198 112154 28250
rect 112206 28198 112258 28250
rect 142718 28198 142770 28250
rect 142822 28198 142874 28250
rect 142926 28198 142978 28250
rect 173438 28198 173490 28250
rect 173542 28198 173594 28250
rect 173646 28198 173698 28250
rect 204158 28198 204210 28250
rect 204262 28198 204314 28250
rect 204366 28198 204418 28250
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 65918 27414 65970 27466
rect 66022 27414 66074 27466
rect 66126 27414 66178 27466
rect 96638 27414 96690 27466
rect 96742 27414 96794 27466
rect 96846 27414 96898 27466
rect 127358 27414 127410 27466
rect 127462 27414 127514 27466
rect 127566 27414 127618 27466
rect 158078 27414 158130 27466
rect 158182 27414 158234 27466
rect 158286 27414 158338 27466
rect 188798 27414 188850 27466
rect 188902 27414 188954 27466
rect 189006 27414 189058 27466
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 50558 26630 50610 26682
rect 50662 26630 50714 26682
rect 50766 26630 50818 26682
rect 81278 26630 81330 26682
rect 81382 26630 81434 26682
rect 81486 26630 81538 26682
rect 111998 26630 112050 26682
rect 112102 26630 112154 26682
rect 112206 26630 112258 26682
rect 142718 26630 142770 26682
rect 142822 26630 142874 26682
rect 142926 26630 142978 26682
rect 173438 26630 173490 26682
rect 173542 26630 173594 26682
rect 173646 26630 173698 26682
rect 204158 26630 204210 26682
rect 204262 26630 204314 26682
rect 204366 26630 204418 26682
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 65918 25846 65970 25898
rect 66022 25846 66074 25898
rect 66126 25846 66178 25898
rect 96638 25846 96690 25898
rect 96742 25846 96794 25898
rect 96846 25846 96898 25898
rect 127358 25846 127410 25898
rect 127462 25846 127514 25898
rect 127566 25846 127618 25898
rect 158078 25846 158130 25898
rect 158182 25846 158234 25898
rect 158286 25846 158338 25898
rect 188798 25846 188850 25898
rect 188902 25846 188954 25898
rect 189006 25846 189058 25898
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 50558 25062 50610 25114
rect 50662 25062 50714 25114
rect 50766 25062 50818 25114
rect 81278 25062 81330 25114
rect 81382 25062 81434 25114
rect 81486 25062 81538 25114
rect 111998 25062 112050 25114
rect 112102 25062 112154 25114
rect 112206 25062 112258 25114
rect 142718 25062 142770 25114
rect 142822 25062 142874 25114
rect 142926 25062 142978 25114
rect 173438 25062 173490 25114
rect 173542 25062 173594 25114
rect 173646 25062 173698 25114
rect 204158 25062 204210 25114
rect 204262 25062 204314 25114
rect 204366 25062 204418 25114
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 65918 24278 65970 24330
rect 66022 24278 66074 24330
rect 66126 24278 66178 24330
rect 96638 24278 96690 24330
rect 96742 24278 96794 24330
rect 96846 24278 96898 24330
rect 127358 24278 127410 24330
rect 127462 24278 127514 24330
rect 127566 24278 127618 24330
rect 158078 24278 158130 24330
rect 158182 24278 158234 24330
rect 158286 24278 158338 24330
rect 188798 24278 188850 24330
rect 188902 24278 188954 24330
rect 189006 24278 189058 24330
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 50558 23494 50610 23546
rect 50662 23494 50714 23546
rect 50766 23494 50818 23546
rect 81278 23494 81330 23546
rect 81382 23494 81434 23546
rect 81486 23494 81538 23546
rect 111998 23494 112050 23546
rect 112102 23494 112154 23546
rect 112206 23494 112258 23546
rect 142718 23494 142770 23546
rect 142822 23494 142874 23546
rect 142926 23494 142978 23546
rect 173438 23494 173490 23546
rect 173542 23494 173594 23546
rect 173646 23494 173698 23546
rect 204158 23494 204210 23546
rect 204262 23494 204314 23546
rect 204366 23494 204418 23546
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 65918 22710 65970 22762
rect 66022 22710 66074 22762
rect 66126 22710 66178 22762
rect 96638 22710 96690 22762
rect 96742 22710 96794 22762
rect 96846 22710 96898 22762
rect 127358 22710 127410 22762
rect 127462 22710 127514 22762
rect 127566 22710 127618 22762
rect 158078 22710 158130 22762
rect 158182 22710 158234 22762
rect 158286 22710 158338 22762
rect 188798 22710 188850 22762
rect 188902 22710 188954 22762
rect 189006 22710 189058 22762
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 50558 21926 50610 21978
rect 50662 21926 50714 21978
rect 50766 21926 50818 21978
rect 81278 21926 81330 21978
rect 81382 21926 81434 21978
rect 81486 21926 81538 21978
rect 111998 21926 112050 21978
rect 112102 21926 112154 21978
rect 112206 21926 112258 21978
rect 142718 21926 142770 21978
rect 142822 21926 142874 21978
rect 142926 21926 142978 21978
rect 173438 21926 173490 21978
rect 173542 21926 173594 21978
rect 173646 21926 173698 21978
rect 204158 21926 204210 21978
rect 204262 21926 204314 21978
rect 204366 21926 204418 21978
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 65918 21142 65970 21194
rect 66022 21142 66074 21194
rect 66126 21142 66178 21194
rect 96638 21142 96690 21194
rect 96742 21142 96794 21194
rect 96846 21142 96898 21194
rect 127358 21142 127410 21194
rect 127462 21142 127514 21194
rect 127566 21142 127618 21194
rect 158078 21142 158130 21194
rect 158182 21142 158234 21194
rect 158286 21142 158338 21194
rect 188798 21142 188850 21194
rect 188902 21142 188954 21194
rect 189006 21142 189058 21194
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 50558 20358 50610 20410
rect 50662 20358 50714 20410
rect 50766 20358 50818 20410
rect 81278 20358 81330 20410
rect 81382 20358 81434 20410
rect 81486 20358 81538 20410
rect 111998 20358 112050 20410
rect 112102 20358 112154 20410
rect 112206 20358 112258 20410
rect 142718 20358 142770 20410
rect 142822 20358 142874 20410
rect 142926 20358 142978 20410
rect 173438 20358 173490 20410
rect 173542 20358 173594 20410
rect 173646 20358 173698 20410
rect 204158 20358 204210 20410
rect 204262 20358 204314 20410
rect 204366 20358 204418 20410
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 65918 19574 65970 19626
rect 66022 19574 66074 19626
rect 66126 19574 66178 19626
rect 96638 19574 96690 19626
rect 96742 19574 96794 19626
rect 96846 19574 96898 19626
rect 127358 19574 127410 19626
rect 127462 19574 127514 19626
rect 127566 19574 127618 19626
rect 158078 19574 158130 19626
rect 158182 19574 158234 19626
rect 158286 19574 158338 19626
rect 188798 19574 188850 19626
rect 188902 19574 188954 19626
rect 189006 19574 189058 19626
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 50558 18790 50610 18842
rect 50662 18790 50714 18842
rect 50766 18790 50818 18842
rect 81278 18790 81330 18842
rect 81382 18790 81434 18842
rect 81486 18790 81538 18842
rect 111998 18790 112050 18842
rect 112102 18790 112154 18842
rect 112206 18790 112258 18842
rect 142718 18790 142770 18842
rect 142822 18790 142874 18842
rect 142926 18790 142978 18842
rect 173438 18790 173490 18842
rect 173542 18790 173594 18842
rect 173646 18790 173698 18842
rect 204158 18790 204210 18842
rect 204262 18790 204314 18842
rect 204366 18790 204418 18842
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 65918 18006 65970 18058
rect 66022 18006 66074 18058
rect 66126 18006 66178 18058
rect 96638 18006 96690 18058
rect 96742 18006 96794 18058
rect 96846 18006 96898 18058
rect 127358 18006 127410 18058
rect 127462 18006 127514 18058
rect 127566 18006 127618 18058
rect 158078 18006 158130 18058
rect 158182 18006 158234 18058
rect 158286 18006 158338 18058
rect 188798 18006 188850 18058
rect 188902 18006 188954 18058
rect 189006 18006 189058 18058
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 50558 17222 50610 17274
rect 50662 17222 50714 17274
rect 50766 17222 50818 17274
rect 81278 17222 81330 17274
rect 81382 17222 81434 17274
rect 81486 17222 81538 17274
rect 111998 17222 112050 17274
rect 112102 17222 112154 17274
rect 112206 17222 112258 17274
rect 142718 17222 142770 17274
rect 142822 17222 142874 17274
rect 142926 17222 142978 17274
rect 173438 17222 173490 17274
rect 173542 17222 173594 17274
rect 173646 17222 173698 17274
rect 204158 17222 204210 17274
rect 204262 17222 204314 17274
rect 204366 17222 204418 17274
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 65918 16438 65970 16490
rect 66022 16438 66074 16490
rect 66126 16438 66178 16490
rect 96638 16438 96690 16490
rect 96742 16438 96794 16490
rect 96846 16438 96898 16490
rect 127358 16438 127410 16490
rect 127462 16438 127514 16490
rect 127566 16438 127618 16490
rect 158078 16438 158130 16490
rect 158182 16438 158234 16490
rect 158286 16438 158338 16490
rect 188798 16438 188850 16490
rect 188902 16438 188954 16490
rect 189006 16438 189058 16490
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 50558 15654 50610 15706
rect 50662 15654 50714 15706
rect 50766 15654 50818 15706
rect 81278 15654 81330 15706
rect 81382 15654 81434 15706
rect 81486 15654 81538 15706
rect 111998 15654 112050 15706
rect 112102 15654 112154 15706
rect 112206 15654 112258 15706
rect 142718 15654 142770 15706
rect 142822 15654 142874 15706
rect 142926 15654 142978 15706
rect 173438 15654 173490 15706
rect 173542 15654 173594 15706
rect 173646 15654 173698 15706
rect 204158 15654 204210 15706
rect 204262 15654 204314 15706
rect 204366 15654 204418 15706
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 65918 14870 65970 14922
rect 66022 14870 66074 14922
rect 66126 14870 66178 14922
rect 96638 14870 96690 14922
rect 96742 14870 96794 14922
rect 96846 14870 96898 14922
rect 127358 14870 127410 14922
rect 127462 14870 127514 14922
rect 127566 14870 127618 14922
rect 158078 14870 158130 14922
rect 158182 14870 158234 14922
rect 158286 14870 158338 14922
rect 188798 14870 188850 14922
rect 188902 14870 188954 14922
rect 189006 14870 189058 14922
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 50558 14086 50610 14138
rect 50662 14086 50714 14138
rect 50766 14086 50818 14138
rect 81278 14086 81330 14138
rect 81382 14086 81434 14138
rect 81486 14086 81538 14138
rect 111998 14086 112050 14138
rect 112102 14086 112154 14138
rect 112206 14086 112258 14138
rect 142718 14086 142770 14138
rect 142822 14086 142874 14138
rect 142926 14086 142978 14138
rect 173438 14086 173490 14138
rect 173542 14086 173594 14138
rect 173646 14086 173698 14138
rect 204158 14086 204210 14138
rect 204262 14086 204314 14138
rect 204366 14086 204418 14138
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 65918 13302 65970 13354
rect 66022 13302 66074 13354
rect 66126 13302 66178 13354
rect 96638 13302 96690 13354
rect 96742 13302 96794 13354
rect 96846 13302 96898 13354
rect 127358 13302 127410 13354
rect 127462 13302 127514 13354
rect 127566 13302 127618 13354
rect 158078 13302 158130 13354
rect 158182 13302 158234 13354
rect 158286 13302 158338 13354
rect 188798 13302 188850 13354
rect 188902 13302 188954 13354
rect 189006 13302 189058 13354
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 50558 12518 50610 12570
rect 50662 12518 50714 12570
rect 50766 12518 50818 12570
rect 81278 12518 81330 12570
rect 81382 12518 81434 12570
rect 81486 12518 81538 12570
rect 111998 12518 112050 12570
rect 112102 12518 112154 12570
rect 112206 12518 112258 12570
rect 142718 12518 142770 12570
rect 142822 12518 142874 12570
rect 142926 12518 142978 12570
rect 173438 12518 173490 12570
rect 173542 12518 173594 12570
rect 173646 12518 173698 12570
rect 204158 12518 204210 12570
rect 204262 12518 204314 12570
rect 204366 12518 204418 12570
rect 156494 12126 156546 12178
rect 156046 12014 156098 12066
rect 163326 12014 163378 12066
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 65918 11734 65970 11786
rect 66022 11734 66074 11786
rect 66126 11734 66178 11786
rect 96638 11734 96690 11786
rect 96742 11734 96794 11786
rect 96846 11734 96898 11786
rect 127358 11734 127410 11786
rect 127462 11734 127514 11786
rect 127566 11734 127618 11786
rect 158078 11734 158130 11786
rect 158182 11734 158234 11786
rect 158286 11734 158338 11786
rect 188798 11734 188850 11786
rect 188902 11734 188954 11786
rect 189006 11734 189058 11786
rect 156606 11566 156658 11618
rect 162542 11566 162594 11618
rect 146862 11454 146914 11506
rect 147310 11454 147362 11506
rect 149214 11454 149266 11506
rect 150446 11454 150498 11506
rect 155262 11454 155314 11506
rect 157726 11454 157778 11506
rect 164670 11454 164722 11506
rect 147534 11342 147586 11394
rect 148206 11342 148258 11394
rect 148766 11342 148818 11394
rect 155598 11342 155650 11394
rect 156718 11342 156770 11394
rect 157166 11342 157218 11394
rect 162430 11342 162482 11394
rect 163102 11342 163154 11394
rect 163998 11342 164050 11394
rect 150110 11230 150162 11282
rect 156494 11230 156546 11282
rect 163438 11230 163490 11282
rect 146190 11118 146242 11170
rect 147870 11118 147922 11170
rect 156942 11118 156994 11170
rect 162654 11118 162706 11170
rect 162878 11118 162930 11170
rect 163326 11118 163378 11170
rect 163662 11118 163714 11170
rect 163886 11118 163938 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 50558 10950 50610 11002
rect 50662 10950 50714 11002
rect 50766 10950 50818 11002
rect 81278 10950 81330 11002
rect 81382 10950 81434 11002
rect 81486 10950 81538 11002
rect 111998 10950 112050 11002
rect 112102 10950 112154 11002
rect 112206 10950 112258 11002
rect 142718 10950 142770 11002
rect 142822 10950 142874 11002
rect 142926 10950 142978 11002
rect 173438 10950 173490 11002
rect 173542 10950 173594 11002
rect 173646 10950 173698 11002
rect 204158 10950 204210 11002
rect 204262 10950 204314 11002
rect 204366 10950 204418 11002
rect 147870 10782 147922 10834
rect 161534 10782 161586 10834
rect 162318 10782 162370 10834
rect 162990 10782 163042 10834
rect 163550 10782 163602 10834
rect 163774 10782 163826 10834
rect 164446 10782 164498 10834
rect 154926 10670 154978 10722
rect 156158 10670 156210 10722
rect 160526 10670 160578 10722
rect 160750 10670 160802 10722
rect 162094 10670 162146 10722
rect 163998 10670 164050 10722
rect 148206 10558 148258 10610
rect 149214 10558 149266 10610
rect 149662 10558 149714 10610
rect 151230 10558 151282 10610
rect 153134 10558 153186 10610
rect 155710 10558 155762 10610
rect 156046 10558 156098 10610
rect 160078 10558 160130 10610
rect 160302 10558 160354 10610
rect 161198 10558 161250 10610
rect 161982 10558 162034 10610
rect 162542 10558 162594 10610
rect 163326 10558 163378 10610
rect 147534 10446 147586 10498
rect 148766 10446 148818 10498
rect 151790 10446 151842 10498
rect 153582 10446 153634 10498
rect 154590 10446 154642 10498
rect 162654 10446 162706 10498
rect 160190 10334 160242 10386
rect 163438 10334 163490 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 65918 10166 65970 10218
rect 66022 10166 66074 10218
rect 66126 10166 66178 10218
rect 96638 10166 96690 10218
rect 96742 10166 96794 10218
rect 96846 10166 96898 10218
rect 127358 10166 127410 10218
rect 127462 10166 127514 10218
rect 127566 10166 127618 10218
rect 158078 10166 158130 10218
rect 158182 10166 158234 10218
rect 158286 10166 158338 10218
rect 188798 10166 188850 10218
rect 188902 10166 188954 10218
rect 189006 10166 189058 10218
rect 139806 9998 139858 10050
rect 140366 9998 140418 10050
rect 139134 9886 139186 9938
rect 139806 9886 139858 9938
rect 140366 9886 140418 9938
rect 148206 9886 148258 9938
rect 157950 9886 158002 9938
rect 161086 9886 161138 9938
rect 140702 9774 140754 9826
rect 148542 9774 148594 9826
rect 149774 9774 149826 9826
rect 151566 9774 151618 9826
rect 151902 9774 151954 9826
rect 152462 9774 152514 9826
rect 154814 9774 154866 9826
rect 155598 9774 155650 9826
rect 155934 9774 155986 9826
rect 156158 9774 156210 9826
rect 156830 9774 156882 9826
rect 157502 9774 157554 9826
rect 150558 9662 150610 9714
rect 155150 9662 155202 9714
rect 157054 9662 157106 9714
rect 161534 9662 161586 9714
rect 161870 9662 161922 9714
rect 141486 9550 141538 9602
rect 148654 9550 148706 9602
rect 149998 9550 150050 9602
rect 154030 9550 154082 9602
rect 155710 9550 155762 9602
rect 156270 9550 156322 9602
rect 156718 9550 156770 9602
rect 157278 9550 157330 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 50558 9382 50610 9434
rect 50662 9382 50714 9434
rect 50766 9382 50818 9434
rect 81278 9382 81330 9434
rect 81382 9382 81434 9434
rect 81486 9382 81538 9434
rect 111998 9382 112050 9434
rect 112102 9382 112154 9434
rect 112206 9382 112258 9434
rect 142718 9382 142770 9434
rect 142822 9382 142874 9434
rect 142926 9382 142978 9434
rect 173438 9382 173490 9434
rect 173542 9382 173594 9434
rect 173646 9382 173698 9434
rect 204158 9382 204210 9434
rect 204262 9382 204314 9434
rect 204366 9382 204418 9434
rect 138686 9214 138738 9266
rect 139582 9214 139634 9266
rect 148430 9214 148482 9266
rect 150110 9214 150162 9266
rect 151566 9214 151618 9266
rect 156046 9214 156098 9266
rect 157166 9214 157218 9266
rect 135326 9102 135378 9154
rect 135998 9102 136050 9154
rect 138238 9102 138290 9154
rect 140254 9102 140306 9154
rect 140926 9102 140978 9154
rect 148542 9102 148594 9154
rect 151006 9102 151058 9154
rect 153358 9102 153410 9154
rect 134542 8990 134594 9042
rect 135550 8990 135602 9042
rect 137678 8990 137730 9042
rect 140814 8990 140866 9042
rect 149326 8990 149378 9042
rect 149550 8990 149602 9042
rect 150670 8990 150722 9042
rect 152126 8990 152178 9042
rect 153918 8990 153970 9042
rect 139134 8878 139186 8930
rect 149662 8878 149714 8930
rect 156494 8878 156546 8930
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 65918 8598 65970 8650
rect 66022 8598 66074 8650
rect 66126 8598 66178 8650
rect 96638 8598 96690 8650
rect 96742 8598 96794 8650
rect 96846 8598 96898 8650
rect 127358 8598 127410 8650
rect 127462 8598 127514 8650
rect 127566 8598 127618 8650
rect 158078 8598 158130 8650
rect 158182 8598 158234 8650
rect 158286 8598 158338 8650
rect 188798 8598 188850 8650
rect 188902 8598 188954 8650
rect 189006 8598 189058 8650
rect 153022 8430 153074 8482
rect 132862 8318 132914 8370
rect 144734 8318 144786 8370
rect 147870 8318 147922 8370
rect 148542 8318 148594 8370
rect 148766 8318 148818 8370
rect 149886 8318 149938 8370
rect 152798 8318 152850 8370
rect 153582 8318 153634 8370
rect 153694 8318 153746 8370
rect 133086 8206 133138 8258
rect 135550 8206 135602 8258
rect 139470 8206 139522 8258
rect 140926 8206 140978 8258
rect 150222 8206 150274 8258
rect 152350 8206 152402 8258
rect 162430 8206 162482 8258
rect 133198 8094 133250 8146
rect 135774 8094 135826 8146
rect 139582 8094 139634 8146
rect 142158 8094 142210 8146
rect 150670 8094 150722 8146
rect 136334 7982 136386 8034
rect 138462 7982 138514 8034
rect 140142 7982 140194 8034
rect 143278 7982 143330 8034
rect 144062 7982 144114 8034
rect 145182 7982 145234 8034
rect 148206 7982 148258 8034
rect 150222 7982 150274 8034
rect 152014 7982 152066 8034
rect 153358 7982 153410 8034
rect 154702 7982 154754 8034
rect 162766 7982 162818 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 50558 7814 50610 7866
rect 50662 7814 50714 7866
rect 50766 7814 50818 7866
rect 81278 7814 81330 7866
rect 81382 7814 81434 7866
rect 81486 7814 81538 7866
rect 111998 7814 112050 7866
rect 112102 7814 112154 7866
rect 112206 7814 112258 7866
rect 142718 7814 142770 7866
rect 142822 7814 142874 7866
rect 142926 7814 142978 7866
rect 173438 7814 173490 7866
rect 173542 7814 173594 7866
rect 173646 7814 173698 7866
rect 204158 7814 204210 7866
rect 204262 7814 204314 7866
rect 204366 7814 204418 7866
rect 132750 7646 132802 7698
rect 136222 7646 136274 7698
rect 140030 7646 140082 7698
rect 147870 7646 147922 7698
rect 151902 7646 151954 7698
rect 153134 7646 153186 7698
rect 153806 7646 153858 7698
rect 160638 7646 160690 7698
rect 132526 7534 132578 7586
rect 133982 7534 134034 7586
rect 135662 7534 135714 7586
rect 138238 7534 138290 7586
rect 139470 7534 139522 7586
rect 142942 7534 142994 7586
rect 148094 7534 148146 7586
rect 151342 7534 151394 7586
rect 151678 7534 151730 7586
rect 152686 7534 152738 7586
rect 161758 7534 161810 7586
rect 162766 7534 162818 7586
rect 163550 7534 163602 7586
rect 131742 7422 131794 7474
rect 134206 7422 134258 7474
rect 135550 7422 135602 7474
rect 137678 7422 137730 7474
rect 139134 7422 139186 7474
rect 140590 7422 140642 7474
rect 141822 7422 141874 7474
rect 144062 7422 144114 7474
rect 145742 7422 145794 7474
rect 146078 7422 146130 7474
rect 146414 7422 146466 7474
rect 147646 7422 147698 7474
rect 149326 7422 149378 7474
rect 150782 7422 150834 7474
rect 150894 7422 150946 7474
rect 151118 7422 151170 7474
rect 152126 7422 152178 7474
rect 152350 7422 152402 7474
rect 152910 7422 152962 7474
rect 153246 7422 153298 7474
rect 161422 7422 161474 7474
rect 162206 7422 162258 7474
rect 162542 7422 162594 7474
rect 162990 7422 163042 7474
rect 163326 7422 163378 7474
rect 150110 7310 150162 7362
rect 151454 7310 151506 7362
rect 152462 7310 152514 7362
rect 154254 7310 154306 7362
rect 154814 7310 154866 7362
rect 155150 7310 155202 7362
rect 161086 7310 161138 7362
rect 164110 7310 164162 7362
rect 152798 7198 152850 7250
rect 162878 7198 162930 7250
rect 163662 7198 163714 7250
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 65918 7030 65970 7082
rect 66022 7030 66074 7082
rect 66126 7030 66178 7082
rect 96638 7030 96690 7082
rect 96742 7030 96794 7082
rect 96846 7030 96898 7082
rect 127358 7030 127410 7082
rect 127462 7030 127514 7082
rect 127566 7030 127618 7082
rect 158078 7030 158130 7082
rect 158182 7030 158234 7082
rect 158286 7030 158338 7082
rect 188798 7030 188850 7082
rect 188902 7030 188954 7082
rect 189006 7030 189058 7082
rect 151902 6750 151954 6802
rect 155374 6750 155426 6802
rect 160638 6750 160690 6802
rect 161534 6750 161586 6802
rect 162766 6750 162818 6802
rect 133086 6638 133138 6690
rect 135214 6638 135266 6690
rect 136334 6638 136386 6690
rect 137230 6638 137282 6690
rect 138238 6638 138290 6690
rect 139022 6638 139074 6690
rect 141822 6638 141874 6690
rect 142494 6638 142546 6690
rect 142942 6638 142994 6690
rect 145406 6638 145458 6690
rect 145854 6638 145906 6690
rect 147646 6638 147698 6690
rect 147982 6638 148034 6690
rect 148654 6638 148706 6690
rect 149998 6638 150050 6690
rect 150334 6638 150386 6690
rect 151118 6638 151170 6690
rect 153358 6638 153410 6690
rect 155598 6638 155650 6690
rect 155822 6638 155874 6690
rect 160974 6638 161026 6690
rect 162654 6638 162706 6690
rect 163886 6638 163938 6690
rect 164334 6638 164386 6690
rect 133198 6526 133250 6578
rect 135774 6526 135826 6578
rect 140366 6526 140418 6578
rect 140702 6526 140754 6578
rect 144622 6526 144674 6578
rect 152126 6526 152178 6578
rect 156606 6526 156658 6578
rect 160302 6526 160354 6578
rect 161422 6526 161474 6578
rect 162878 6526 162930 6578
rect 134654 6414 134706 6466
rect 137902 6414 137954 6466
rect 138910 6414 138962 6466
rect 144286 6414 144338 6466
rect 147310 6414 147362 6466
rect 148318 6414 148370 6466
rect 154030 6414 154082 6466
rect 159966 6414 160018 6466
rect 160526 6414 160578 6466
rect 160750 6414 160802 6466
rect 161646 6414 161698 6466
rect 163102 6414 163154 6466
rect 163774 6414 163826 6466
rect 164446 6414 164498 6466
rect 164558 6414 164610 6466
rect 165118 6414 165170 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 50558 6246 50610 6298
rect 50662 6246 50714 6298
rect 50766 6246 50818 6298
rect 81278 6246 81330 6298
rect 81382 6246 81434 6298
rect 81486 6246 81538 6298
rect 111998 6246 112050 6298
rect 112102 6246 112154 6298
rect 112206 6246 112258 6298
rect 142718 6246 142770 6298
rect 142822 6246 142874 6298
rect 142926 6246 142978 6298
rect 173438 6246 173490 6298
rect 173542 6246 173594 6298
rect 173646 6246 173698 6298
rect 204158 6246 204210 6298
rect 204262 6246 204314 6298
rect 204366 6246 204418 6298
rect 135550 6078 135602 6130
rect 138014 6078 138066 6130
rect 145294 6078 145346 6130
rect 149662 6078 149714 6130
rect 156830 6078 156882 6130
rect 157950 6078 158002 6130
rect 159294 6078 159346 6130
rect 159630 6078 159682 6130
rect 159854 6078 159906 6130
rect 161198 6078 161250 6130
rect 162318 6078 162370 6130
rect 164894 6078 164946 6130
rect 137230 5966 137282 6018
rect 139806 5966 139858 6018
rect 145070 5966 145122 6018
rect 149886 5966 149938 6018
rect 151454 5966 151506 6018
rect 152686 5966 152738 6018
rect 154702 5966 154754 6018
rect 160414 5966 160466 6018
rect 160638 5966 160690 6018
rect 162990 5966 163042 6018
rect 163214 5966 163266 6018
rect 163998 5966 164050 6018
rect 136446 5854 136498 5906
rect 138910 5854 138962 5906
rect 139134 5854 139186 5906
rect 140142 5854 140194 5906
rect 141822 5854 141874 5906
rect 143950 5854 144002 5906
rect 146078 5854 146130 5906
rect 146750 5854 146802 5906
rect 147198 5854 147250 5906
rect 148542 5854 148594 5906
rect 149438 5854 149490 5906
rect 150110 5854 150162 5906
rect 151342 5854 151394 5906
rect 152126 5854 152178 5906
rect 152462 5854 152514 5906
rect 153918 5854 153970 5906
rect 154142 5854 154194 5906
rect 156382 5854 156434 5906
rect 160190 5854 160242 5906
rect 160750 5854 160802 5906
rect 161758 5854 161810 5906
rect 162542 5854 162594 5906
rect 163326 5854 163378 5906
rect 163550 5854 163602 5906
rect 164110 5854 164162 5906
rect 164222 5854 164274 5906
rect 164446 5854 164498 5906
rect 165118 5854 165170 5906
rect 165566 5854 165618 5906
rect 135102 5742 135154 5794
rect 139470 5742 139522 5794
rect 140590 5742 140642 5794
rect 141262 5742 141314 5794
rect 149102 5742 149154 5794
rect 150222 5742 150274 5794
rect 150782 5742 150834 5794
rect 155934 5742 155986 5794
rect 157390 5742 157442 5794
rect 165006 5742 165058 5794
rect 153134 5630 153186 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 65918 5462 65970 5514
rect 66022 5462 66074 5514
rect 66126 5462 66178 5514
rect 96638 5462 96690 5514
rect 96742 5462 96794 5514
rect 96846 5462 96898 5514
rect 127358 5462 127410 5514
rect 127462 5462 127514 5514
rect 127566 5462 127618 5514
rect 158078 5462 158130 5514
rect 158182 5462 158234 5514
rect 158286 5462 158338 5514
rect 188798 5462 188850 5514
rect 188902 5462 188954 5514
rect 189006 5462 189058 5514
rect 130510 5294 130562 5346
rect 131294 5294 131346 5346
rect 131742 5294 131794 5346
rect 133758 5294 133810 5346
rect 134206 5294 134258 5346
rect 134542 5294 134594 5346
rect 135774 5294 135826 5346
rect 152574 5294 152626 5346
rect 153022 5294 153074 5346
rect 155150 5294 155202 5346
rect 156382 5294 156434 5346
rect 6414 5182 6466 5234
rect 49758 5182 49810 5234
rect 52110 5182 52162 5234
rect 55134 5182 55186 5234
rect 57822 5182 57874 5234
rect 59950 5182 60002 5234
rect 63198 5182 63250 5234
rect 65886 5182 65938 5234
rect 68574 5182 68626 5234
rect 92766 5182 92818 5234
rect 93774 5182 93826 5234
rect 97470 5182 97522 5234
rect 98366 5182 98418 5234
rect 102062 5182 102114 5234
rect 105534 5182 105586 5234
rect 106542 5182 106594 5234
rect 109230 5182 109282 5234
rect 110350 5182 110402 5234
rect 110798 5182 110850 5234
rect 113374 5182 113426 5234
rect 114382 5182 114434 5234
rect 117630 5182 117682 5234
rect 118526 5182 118578 5234
rect 121214 5182 121266 5234
rect 122222 5182 122274 5234
rect 125582 5182 125634 5234
rect 126590 5182 126642 5234
rect 130062 5182 130114 5234
rect 130398 5182 130450 5234
rect 132078 5182 132130 5234
rect 132638 5182 132690 5234
rect 133422 5182 133474 5234
rect 137454 5182 137506 5234
rect 145406 5182 145458 5234
rect 145854 5182 145906 5234
rect 157950 5182 158002 5234
rect 161870 5182 161922 5234
rect 162878 5182 162930 5234
rect 5966 5070 6018 5122
rect 50094 5070 50146 5122
rect 52782 5070 52834 5122
rect 55470 5070 55522 5122
rect 58158 5070 58210 5122
rect 60846 5070 60898 5122
rect 63534 5070 63586 5122
rect 66222 5070 66274 5122
rect 68910 5070 68962 5122
rect 93326 5070 93378 5122
rect 97918 5070 97970 5122
rect 101614 5070 101666 5122
rect 106094 5070 106146 5122
rect 109678 5070 109730 5122
rect 110014 5070 110066 5122
rect 113934 5070 113986 5122
rect 118078 5070 118130 5122
rect 121774 5070 121826 5122
rect 126142 5070 126194 5122
rect 131182 5070 131234 5122
rect 133646 5070 133698 5122
rect 135326 5070 135378 5122
rect 136894 5070 136946 5122
rect 138126 5070 138178 5122
rect 138910 5070 138962 5122
rect 141822 5070 141874 5122
rect 142494 5070 142546 5122
rect 143054 5070 143106 5122
rect 144286 5070 144338 5122
rect 144958 5070 145010 5122
rect 146750 5070 146802 5122
rect 148990 5070 149042 5122
rect 150334 5070 150386 5122
rect 150558 5070 150610 5122
rect 152014 5070 152066 5122
rect 152238 5070 152290 5122
rect 152574 5070 152626 5122
rect 153470 5070 153522 5122
rect 153694 5070 153746 5122
rect 154030 5070 154082 5122
rect 154590 5070 154642 5122
rect 155374 5070 155426 5122
rect 155598 5070 155650 5122
rect 155710 5070 155762 5122
rect 156158 5070 156210 5122
rect 156718 5070 156770 5122
rect 157166 5070 157218 5122
rect 157278 5070 157330 5122
rect 157390 5070 157442 5122
rect 157838 5070 157890 5122
rect 160526 5070 160578 5122
rect 161086 5070 161138 5122
rect 161534 5070 161586 5122
rect 162318 5070 162370 5122
rect 162766 5070 162818 5122
rect 163326 5070 163378 5122
rect 163662 5070 163714 5122
rect 163774 5070 163826 5122
rect 163998 5070 164050 5122
rect 164782 5070 164834 5122
rect 165230 5070 165282 5122
rect 165678 5070 165730 5122
rect 166126 5070 166178 5122
rect 166238 5070 166290 5122
rect 101054 4958 101106 5010
rect 131630 4958 131682 5010
rect 132190 4958 132242 5010
rect 134094 4958 134146 5010
rect 135662 4958 135714 5010
rect 137006 4958 137058 5010
rect 138014 4958 138066 5010
rect 140366 4958 140418 5010
rect 140702 4958 140754 5010
rect 148206 4958 148258 5010
rect 148542 4958 148594 5010
rect 152462 4958 152514 5010
rect 153918 4958 153970 5010
rect 158286 4958 158338 5010
rect 160302 4958 160354 5010
rect 161758 4958 161810 5010
rect 162990 4958 163042 5010
rect 5630 4846 5682 4898
rect 50430 4846 50482 4898
rect 53118 4846 53170 4898
rect 55806 4846 55858 4898
rect 58494 4846 58546 4898
rect 61182 4846 61234 4898
rect 63870 4846 63922 4898
rect 66558 4846 66610 4898
rect 69246 4846 69298 4898
rect 136446 4846 136498 4898
rect 140814 4846 140866 4898
rect 146862 4846 146914 4898
rect 154814 4846 154866 4898
rect 155038 4846 155090 4898
rect 156494 4846 156546 4898
rect 158062 4846 158114 4898
rect 160862 4846 160914 4898
rect 164446 4846 164498 4898
rect 165342 4846 165394 4898
rect 165454 4846 165506 4898
rect 166350 4846 166402 4898
rect 166910 4846 166962 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 50558 4678 50610 4730
rect 50662 4678 50714 4730
rect 50766 4678 50818 4730
rect 81278 4678 81330 4730
rect 81382 4678 81434 4730
rect 81486 4678 81538 4730
rect 111998 4678 112050 4730
rect 112102 4678 112154 4730
rect 112206 4678 112258 4730
rect 142718 4678 142770 4730
rect 142822 4678 142874 4730
rect 142926 4678 142978 4730
rect 173438 4678 173490 4730
rect 173542 4678 173594 4730
rect 173646 4678 173698 4730
rect 204158 4678 204210 4730
rect 204262 4678 204314 4730
rect 204366 4678 204418 4730
rect 33182 4510 33234 4562
rect 35646 4510 35698 4562
rect 44494 4510 44546 4562
rect 46958 4510 47010 4562
rect 88062 4510 88114 4562
rect 88958 4510 89010 4562
rect 139246 4510 139298 4562
rect 145182 4510 145234 4562
rect 149102 4510 149154 4562
rect 149662 4510 149714 4562
rect 149886 4510 149938 4562
rect 150670 4510 150722 4562
rect 151006 4510 151058 4562
rect 155038 4510 155090 4562
rect 155262 4510 155314 4562
rect 155374 4510 155426 4562
rect 160862 4510 160914 4562
rect 161422 4510 161474 4562
rect 163662 4510 163714 4562
rect 163774 4510 163826 4562
rect 52558 4398 52610 4450
rect 138798 4398 138850 4450
rect 144958 4398 145010 4450
rect 150110 4398 150162 4450
rect 150222 4398 150274 4450
rect 152798 4398 152850 4450
rect 153694 4398 153746 4450
rect 155822 4398 155874 4450
rect 156494 4398 156546 4450
rect 162766 4398 162818 4450
rect 164222 4398 164274 4450
rect 5966 4286 6018 4338
rect 32510 4286 32562 4338
rect 44046 4286 44098 4338
rect 51998 4286 52050 4338
rect 57598 4286 57650 4338
rect 68350 4286 68402 4338
rect 78878 4286 78930 4338
rect 79550 4286 79602 4338
rect 81342 4286 81394 4338
rect 87054 4286 87106 4338
rect 137342 4286 137394 4338
rect 140254 4286 140306 4338
rect 140478 4286 140530 4338
rect 140926 4286 140978 4338
rect 142270 4286 142322 4338
rect 143502 4286 143554 4338
rect 146078 4286 146130 4338
rect 146638 4286 146690 4338
rect 147086 4286 147138 4338
rect 148430 4286 148482 4338
rect 148878 4286 148930 4338
rect 149438 4286 149490 4338
rect 151454 4286 151506 4338
rect 154590 4286 154642 4338
rect 155598 4286 155650 4338
rect 156270 4286 156322 4338
rect 161646 4286 161698 4338
rect 161982 4286 162034 4338
rect 162206 4286 162258 4338
rect 162430 4286 162482 4338
rect 162990 4286 163042 4338
rect 163998 4286 164050 4338
rect 130846 4174 130898 4226
rect 131294 4174 131346 4226
rect 133758 4174 133810 4226
rect 135326 4174 135378 4226
rect 143054 4174 143106 4226
rect 151230 4174 151282 4226
rect 165678 4174 165730 4226
rect 4062 4062 4114 4114
rect 30606 4062 30658 4114
rect 41694 4062 41746 4114
rect 49758 4062 49810 4114
rect 58606 4062 58658 4114
rect 69358 4062 69410 4114
rect 76638 4062 76690 4114
rect 84702 4062 84754 4114
rect 161758 4062 161810 4114
rect 163326 4062 163378 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 65918 3894 65970 3946
rect 66022 3894 66074 3946
rect 66126 3894 66178 3946
rect 96638 3894 96690 3946
rect 96742 3894 96794 3946
rect 96846 3894 96898 3946
rect 127358 3894 127410 3946
rect 127462 3894 127514 3946
rect 127566 3894 127618 3946
rect 158078 3894 158130 3946
rect 158182 3894 158234 3946
rect 158286 3894 158338 3946
rect 188798 3894 188850 3946
rect 188902 3894 188954 3946
rect 189006 3894 189058 3946
rect 147870 3726 147922 3778
rect 148766 3726 148818 3778
rect 161534 3726 161586 3778
rect 162318 3726 162370 3778
rect 28590 3614 28642 3666
rect 31502 3614 31554 3666
rect 33182 3614 33234 3666
rect 36318 3614 36370 3666
rect 39230 3614 39282 3666
rect 42926 3614 42978 3666
rect 44382 3614 44434 3666
rect 47630 3614 47682 3666
rect 50542 3614 50594 3666
rect 52894 3614 52946 3666
rect 56030 3614 56082 3666
rect 60510 3614 60562 3666
rect 63982 3614 64034 3666
rect 67454 3614 67506 3666
rect 74286 3614 74338 3666
rect 77198 3614 77250 3666
rect 78878 3614 78930 3666
rect 82014 3614 82066 3666
rect 142830 3614 142882 3666
rect 147422 3614 147474 3666
rect 147870 3614 147922 3666
rect 148318 3614 148370 3666
rect 150334 3614 150386 3666
rect 152798 3614 152850 3666
rect 154478 3614 154530 3666
rect 156158 3614 156210 3666
rect 162318 3614 162370 3666
rect 211598 3614 211650 3666
rect 213950 3614 214002 3666
rect 216638 3614 216690 3666
rect 30942 3502 30994 3554
rect 35422 3502 35474 3554
rect 38670 3502 38722 3554
rect 42366 3502 42418 3554
rect 46734 3502 46786 3554
rect 49982 3502 50034 3554
rect 51886 3502 51938 3554
rect 55022 3502 55074 3554
rect 59502 3502 59554 3554
rect 62974 3502 63026 3554
rect 66446 3502 66498 3554
rect 70926 3502 70978 3554
rect 76526 3502 76578 3554
rect 81118 3502 81170 3554
rect 84366 3502 84418 3554
rect 88734 3502 88786 3554
rect 148766 3502 148818 3554
rect 150894 3502 150946 3554
rect 151342 3502 151394 3554
rect 152014 3502 152066 3554
rect 152238 3502 152290 3554
rect 152462 3502 152514 3554
rect 152686 3502 152738 3554
rect 153358 3502 153410 3554
rect 154030 3502 154082 3554
rect 155038 3502 155090 3554
rect 155710 3502 155762 3554
rect 162654 3502 162706 3554
rect 165678 3502 165730 3554
rect 170718 3502 170770 3554
rect 176094 3502 176146 3554
rect 178782 3502 178834 3554
rect 184718 3502 184770 3554
rect 186846 3502 186898 3554
rect 189534 3502 189586 3554
rect 192334 3502 192386 3554
rect 197934 3502 197986 3554
rect 205998 3502 206050 3554
rect 40574 3390 40626 3442
rect 84926 3390 84978 3442
rect 86942 3390 86994 3442
rect 89630 3390 89682 3442
rect 89854 3390 89906 3442
rect 90190 3390 90242 3442
rect 92654 3390 92706 3442
rect 93102 3390 93154 3442
rect 93438 3390 93490 3442
rect 95006 3390 95058 3442
rect 95230 3390 95282 3442
rect 95566 3390 95618 3442
rect 97694 3390 97746 3442
rect 97918 3390 97970 3442
rect 98254 3390 98306 3442
rect 100270 3390 100322 3442
rect 100718 3390 100770 3442
rect 101054 3390 101106 3442
rect 103070 3390 103122 3442
rect 103294 3390 103346 3442
rect 103630 3390 103682 3442
rect 105758 3390 105810 3442
rect 105982 3390 106034 3442
rect 106318 3390 106370 3442
rect 107886 3390 107938 3442
rect 108670 3390 108722 3442
rect 109006 3390 109058 3442
rect 111694 3390 111746 3442
rect 112142 3390 112194 3442
rect 112478 3390 112530 3442
rect 113822 3390 113874 3442
rect 114046 3390 114098 3442
rect 114382 3390 114434 3442
rect 116510 3390 116562 3442
rect 116734 3390 116786 3442
rect 117070 3390 117122 3442
rect 119310 3390 119362 3442
rect 119758 3390 119810 3442
rect 120094 3390 120146 3442
rect 121886 3390 121938 3442
rect 122110 3390 122162 3442
rect 124574 3390 124626 3442
rect 124798 3390 124850 3442
rect 125134 3390 125186 3442
rect 126926 3390 126978 3442
rect 127486 3390 127538 3442
rect 127822 3390 127874 3442
rect 129950 3390 130002 3442
rect 130174 3390 130226 3442
rect 130510 3390 130562 3442
rect 132638 3390 132690 3442
rect 132862 3390 132914 3442
rect 133198 3390 133250 3442
rect 135326 3390 135378 3442
rect 135550 3390 135602 3442
rect 135886 3390 135938 3442
rect 138350 3390 138402 3442
rect 138798 3390 138850 3442
rect 139134 3390 139186 3442
rect 140702 3390 140754 3442
rect 140926 3390 140978 3442
rect 141262 3390 141314 3442
rect 143390 3390 143442 3442
rect 143614 3390 143666 3442
rect 143950 3390 144002 3442
rect 145966 3390 146018 3442
rect 146414 3390 146466 3442
rect 146750 3390 146802 3442
rect 148990 3390 149042 3442
rect 149326 3390 149378 3442
rect 153022 3390 153074 3442
rect 155262 3390 155314 3442
rect 156606 3390 156658 3442
rect 157390 3390 157442 3442
rect 157838 3390 157890 3442
rect 158174 3390 158226 3442
rect 159518 3390 159570 3442
rect 160078 3390 160130 3442
rect 161982 3390 162034 3442
rect 162990 3390 163042 3442
rect 163326 3390 163378 3442
rect 163662 3390 163714 3442
rect 165006 3390 165058 3442
rect 165454 3390 165506 3442
rect 167582 3390 167634 3442
rect 168142 3390 168194 3442
rect 170270 3390 170322 3442
rect 172622 3390 172674 3442
rect 173182 3390 173234 3442
rect 173518 3390 173570 3442
rect 175646 3390 175698 3442
rect 178334 3390 178386 3442
rect 181022 3390 181074 3442
rect 181582 3390 181634 3442
rect 184046 3390 184098 3442
rect 186398 3390 186450 3442
rect 189086 3390 189138 3442
rect 191662 3390 191714 3442
rect 194462 3390 194514 3442
rect 195022 3390 195074 3442
rect 197150 3390 197202 3442
rect 197374 3390 197426 3442
rect 199278 3390 199330 3442
rect 200062 3390 200114 3442
rect 200622 3390 200674 3442
rect 203086 3390 203138 3442
rect 203534 3390 203586 3442
rect 204094 3390 204146 3442
rect 205214 3390 205266 3442
rect 205438 3390 205490 3442
rect 207902 3390 207954 3442
rect 208126 3390 208178 3442
rect 208686 3390 208738 3442
rect 210702 3390 210754 3442
rect 211150 3390 211202 3442
rect 213278 3390 213330 3442
rect 213502 3390 213554 3442
rect 215966 3390 216018 3442
rect 216190 3390 216242 3442
rect 6526 3278 6578 3330
rect 9326 3278 9378 3330
rect 11902 3278 11954 3330
rect 14590 3278 14642 3330
rect 17278 3278 17330 3330
rect 19966 3278 20018 3330
rect 22654 3278 22706 3330
rect 25342 3278 25394 3330
rect 71934 3278 71986 3330
rect 122446 3278 122498 3330
rect 159742 3278 159794 3330
rect 167806 3278 167858 3330
rect 170494 3278 170546 3330
rect 175870 3278 175922 3330
rect 178558 3278 178610 3330
rect 181246 3278 181298 3330
rect 184494 3278 184546 3330
rect 186622 3278 186674 3330
rect 189310 3278 189362 3330
rect 192110 3278 192162 3330
rect 194686 3278 194738 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 50558 3110 50610 3162
rect 50662 3110 50714 3162
rect 50766 3110 50818 3162
rect 81278 3110 81330 3162
rect 81382 3110 81434 3162
rect 81486 3110 81538 3162
rect 111998 3110 112050 3162
rect 112102 3110 112154 3162
rect 112206 3110 112258 3162
rect 142718 3110 142770 3162
rect 142822 3110 142874 3162
rect 142926 3110 142978 3162
rect 173438 3110 173490 3162
rect 173542 3110 173594 3162
rect 173646 3110 173698 3162
rect 204158 3110 204210 3162
rect 204262 3110 204314 3162
rect 204366 3110 204418 3162
<< metal2 >>
rect 2912 49200 3024 50000
rect 6944 49200 7056 50000
rect 10976 49200 11088 50000
rect 15008 49200 15120 50000
rect 19040 49200 19152 50000
rect 23072 49200 23184 50000
rect 27104 49200 27216 50000
rect 31136 49200 31248 50000
rect 35168 49200 35280 50000
rect 39200 49200 39312 50000
rect 43232 49200 43344 50000
rect 47264 49200 47376 50000
rect 51296 49200 51408 50000
rect 55328 49200 55440 50000
rect 59360 49200 59472 50000
rect 63392 49200 63504 50000
rect 67424 49200 67536 50000
rect 71456 49200 71568 50000
rect 75488 49200 75600 50000
rect 79520 49200 79632 50000
rect 83552 49200 83664 50000
rect 87584 49200 87696 50000
rect 91616 49200 91728 50000
rect 95648 49200 95760 50000
rect 99680 49200 99792 50000
rect 103712 49200 103824 50000
rect 107744 49200 107856 50000
rect 111776 49200 111888 50000
rect 115808 49200 115920 50000
rect 119840 49200 119952 50000
rect 123872 49200 123984 50000
rect 127904 49200 128016 50000
rect 131936 49200 132048 50000
rect 135968 49200 136080 50000
rect 140000 49200 140112 50000
rect 144032 49200 144144 50000
rect 148064 49200 148176 50000
rect 152096 49200 152208 50000
rect 156128 49200 156240 50000
rect 160160 49200 160272 50000
rect 164192 49200 164304 50000
rect 168224 49200 168336 50000
rect 172256 49200 172368 50000
rect 176288 49200 176400 50000
rect 180320 49200 180432 50000
rect 184352 49200 184464 50000
rect 188384 49200 188496 50000
rect 192416 49200 192528 50000
rect 196448 49200 196560 50000
rect 200480 49200 200592 50000
rect 204512 49200 204624 50000
rect 208544 49200 208656 50000
rect 212576 49200 212688 50000
rect 216608 49200 216720 50000
rect 2940 37156 2996 49200
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 6972 46004 7028 49200
rect 11004 46004 11060 49200
rect 15036 46004 15092 49200
rect 19068 46004 19124 49200
rect 23100 46004 23156 49200
rect 27132 46450 27188 49200
rect 31164 47012 31220 49200
rect 31164 46956 31668 47012
rect 27132 46398 27134 46450
rect 27186 46398 27188 46450
rect 27132 46386 27188 46398
rect 27804 46450 27860 46462
rect 27804 46398 27806 46450
rect 27858 46398 27860 46450
rect 6972 46002 7476 46004
rect 6972 45950 6974 46002
rect 7026 45950 7476 46002
rect 6972 45948 7476 45950
rect 6972 45938 7028 45948
rect 7420 45890 7476 45948
rect 11004 46002 11284 46004
rect 11004 45950 11006 46002
rect 11058 45950 11284 46002
rect 11004 45948 11284 45950
rect 11004 45938 11060 45948
rect 7420 45838 7422 45890
rect 7474 45838 7476 45890
rect 7420 45826 7476 45838
rect 11228 45890 11284 45948
rect 15036 46002 15316 46004
rect 15036 45950 15038 46002
rect 15090 45950 15316 46002
rect 15036 45948 15316 45950
rect 15036 45938 15092 45948
rect 11228 45838 11230 45890
rect 11282 45838 11284 45890
rect 11228 45826 11284 45838
rect 15260 45890 15316 45948
rect 19068 46002 19348 46004
rect 19068 45950 19070 46002
rect 19122 45950 19348 46002
rect 19068 45948 19348 45950
rect 19068 45938 19124 45948
rect 15260 45838 15262 45890
rect 15314 45838 15316 45890
rect 15260 45826 15316 45838
rect 15820 45890 15876 45902
rect 15820 45838 15822 45890
rect 15874 45838 15876 45890
rect 12348 45778 12404 45790
rect 12348 45726 12350 45778
rect 12402 45726 12404 45778
rect 7196 45666 7252 45678
rect 7196 45614 7198 45666
rect 7250 45614 7252 45666
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 2940 37090 2996 37100
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 5964 5236 6020 5246
rect 5964 5122 6020 5180
rect 6412 5236 6468 5246
rect 6412 5142 6468 5180
rect 7196 5236 7252 45614
rect 12348 45108 12404 45726
rect 12348 45042 12404 45052
rect 15820 7588 15876 45838
rect 19292 45890 19348 45948
rect 23100 46002 23380 46004
rect 23100 45950 23102 46002
rect 23154 45950 23380 46002
rect 23100 45948 23380 45950
rect 23100 45938 23156 45948
rect 19292 45838 19294 45890
rect 19346 45838 19348 45890
rect 19292 45826 19348 45838
rect 19852 45892 19908 45902
rect 19852 45798 19908 45836
rect 22652 45892 22708 45902
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 22652 9268 22708 45836
rect 23324 45890 23380 45948
rect 27804 46002 27860 46398
rect 27804 45950 27806 46002
rect 27858 45950 27860 46002
rect 27804 45938 27860 45950
rect 28364 46450 28420 46462
rect 28364 46398 28366 46450
rect 28418 46398 28420 46450
rect 23324 45838 23326 45890
rect 23378 45838 23380 45890
rect 23324 45826 23380 45838
rect 23884 45890 23940 45902
rect 23884 45838 23886 45890
rect 23938 45838 23940 45890
rect 23884 26068 23940 45838
rect 28364 45890 28420 46398
rect 31612 46004 31668 46956
rect 35196 46900 35252 49200
rect 35196 46844 35588 46900
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 31612 45910 31668 45948
rect 32172 46004 32228 46014
rect 28364 45838 28366 45890
rect 28418 45838 28420 45890
rect 28364 45826 28420 45838
rect 28924 45890 28980 45902
rect 28924 45838 28926 45890
rect 28978 45838 28980 45890
rect 23884 26002 23940 26012
rect 28924 12740 28980 45838
rect 32172 45890 32228 45948
rect 35420 46004 35476 46014
rect 35532 46004 35588 46844
rect 39228 46004 39284 49200
rect 35420 46002 36036 46004
rect 35420 45950 35422 46002
rect 35474 45950 36036 46002
rect 35420 45948 36036 45950
rect 35420 45938 35476 45948
rect 32172 45838 32174 45890
rect 32226 45838 32228 45890
rect 32172 45826 32228 45838
rect 32732 45890 32788 45902
rect 32732 45838 32734 45890
rect 32786 45838 32788 45890
rect 32732 45444 32788 45838
rect 35980 45890 36036 45948
rect 39228 46002 39844 46004
rect 39228 45950 39230 46002
rect 39282 45950 39844 46002
rect 39228 45948 39844 45950
rect 39228 45938 39284 45948
rect 35980 45838 35982 45890
rect 36034 45838 36036 45890
rect 35980 45826 36036 45838
rect 36540 45892 36596 45902
rect 36540 45798 36596 45836
rect 37772 45892 37828 45902
rect 32732 45378 32788 45388
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 37772 15988 37828 45836
rect 39788 45890 39844 45948
rect 39788 45838 39790 45890
rect 39842 45838 39844 45890
rect 39788 45826 39844 45838
rect 40236 46002 40292 46014
rect 40236 45950 40238 46002
rect 40290 45950 40292 46002
rect 37772 15922 37828 15932
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 28924 12674 28980 12684
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 40236 11284 40292 45950
rect 43148 46004 43204 46014
rect 43260 46004 43316 49200
rect 47292 47460 47348 49200
rect 47292 47404 47796 47460
rect 47740 46114 47796 47404
rect 51324 46564 51380 49200
rect 55356 47068 55412 49200
rect 59388 47460 59444 49200
rect 59388 47404 59780 47460
rect 55356 47012 55860 47068
rect 51324 46508 51828 46564
rect 47740 46062 47742 46114
rect 47794 46062 47796 46114
rect 47740 46050 47796 46062
rect 51772 46114 51828 46508
rect 51772 46062 51774 46114
rect 51826 46062 51828 46114
rect 51772 46050 51828 46062
rect 55804 46114 55860 47012
rect 55804 46062 55806 46114
rect 55858 46062 55860 46114
rect 55804 46050 55860 46062
rect 59724 46114 59780 47404
rect 59724 46062 59726 46114
rect 59778 46062 59780 46114
rect 59724 46050 59780 46062
rect 63420 46116 63476 49200
rect 65916 46284 66180 46294
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 65916 46218 66180 46228
rect 63532 46116 63588 46126
rect 63420 46114 63588 46116
rect 63420 46062 63534 46114
rect 63586 46062 63588 46114
rect 63420 46060 63588 46062
rect 63532 46050 63588 46060
rect 43148 46002 43652 46004
rect 43148 45950 43150 46002
rect 43202 45950 43652 46002
rect 43148 45948 43652 45950
rect 43148 45938 43204 45948
rect 43596 45890 43652 45948
rect 67452 46002 67508 49200
rect 67452 45950 67454 46002
rect 67506 45950 67508 46002
rect 67452 45938 67508 45950
rect 71484 46002 71540 49200
rect 71484 45950 71486 46002
rect 71538 45950 71540 46002
rect 71484 45938 71540 45950
rect 43596 45838 43598 45890
rect 43650 45838 43652 45890
rect 43596 45826 43652 45838
rect 44156 45892 44212 45902
rect 44156 45798 44212 45836
rect 47852 45892 47908 45902
rect 42812 45444 42868 45454
rect 42812 14308 42868 45388
rect 47852 19348 47908 45836
rect 50092 45890 50148 45902
rect 50092 45838 50094 45890
rect 50146 45838 50148 45890
rect 50092 45668 50148 45838
rect 54124 45892 54180 45902
rect 54124 45798 54180 45836
rect 55132 45892 55188 45902
rect 55132 45798 55188 45836
rect 58044 45892 58100 45902
rect 50092 45602 50148 45612
rect 50540 45668 50596 45706
rect 50540 45602 50596 45612
rect 52892 45668 52948 45678
rect 50556 45500 50820 45510
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50556 45434 50820 45444
rect 50556 43932 50820 43942
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50556 43866 50820 43876
rect 50556 42364 50820 42374
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50556 42298 50820 42308
rect 50556 40796 50820 40806
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50556 40730 50820 40740
rect 50556 39228 50820 39238
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50556 39162 50820 39172
rect 50556 37660 50820 37670
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50556 37594 50820 37604
rect 50556 36092 50820 36102
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50556 36026 50820 36036
rect 50556 34524 50820 34534
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50556 34458 50820 34468
rect 50556 32956 50820 32966
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50556 32890 50820 32900
rect 50556 31388 50820 31398
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50556 31322 50820 31332
rect 50556 29820 50820 29830
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50556 29754 50820 29764
rect 50556 28252 50820 28262
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50556 28186 50820 28196
rect 50556 26684 50820 26694
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50556 26618 50820 26628
rect 50556 25116 50820 25126
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50556 25050 50820 25060
rect 50556 23548 50820 23558
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50556 23482 50820 23492
rect 50556 21980 50820 21990
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50556 21914 50820 21924
rect 50556 20412 50820 20422
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50556 20346 50820 20356
rect 47852 19282 47908 19292
rect 50556 18844 50820 18854
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50556 18778 50820 18788
rect 50556 17276 50820 17286
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50556 17210 50820 17220
rect 50556 15708 50820 15718
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50556 15642 50820 15652
rect 42812 14242 42868 14252
rect 50556 14140 50820 14150
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50556 14074 50820 14084
rect 50556 12572 50820 12582
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50556 12506 50820 12516
rect 40236 11218 40292 11228
rect 52892 11172 52948 45612
rect 52892 11106 52948 11116
rect 55132 26068 55188 26078
rect 50556 11004 50820 11014
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50556 10938 50820 10948
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 50556 9436 50820 9446
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50556 9370 50820 9380
rect 22652 9202 22708 9212
rect 52108 9268 52164 9278
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 50556 7868 50820 7878
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50556 7802 50820 7812
rect 15820 7522 15876 7532
rect 49756 7588 49812 7598
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 33180 6916 33236 6926
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 7196 5170 7252 5180
rect 31500 5796 31556 5806
rect 5964 5070 5966 5122
rect 6018 5070 6020 5122
rect 5964 5058 6020 5070
rect 5628 4898 5684 4910
rect 5628 4846 5630 4898
rect 5682 4846 5684 4898
rect 5628 4340 5684 4846
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 5964 4340 6020 4350
rect 5628 4338 6020 4340
rect 5628 4286 5966 4338
rect 6018 4286 6020 4338
rect 5628 4284 6020 4286
rect 5964 4274 6020 4284
rect 4060 4116 4116 4126
rect 3612 4114 4116 4116
rect 3612 4062 4062 4114
rect 4114 4062 4116 4114
rect 3612 4060 4116 4062
rect 3612 800 3668 4060
rect 4060 4050 4116 4060
rect 30604 4114 30660 4126
rect 30604 4062 30606 4114
rect 30658 4062 30660 4114
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 27804 3668 27860 3678
rect 6524 3332 6580 3342
rect 9324 3332 9380 3342
rect 11900 3332 11956 3342
rect 14588 3332 14644 3342
rect 17276 3332 17332 3342
rect 19964 3332 20020 3342
rect 22652 3332 22708 3342
rect 25340 3332 25396 3342
rect 6300 3330 6580 3332
rect 6300 3278 6526 3330
rect 6578 3278 6580 3330
rect 6300 3276 6580 3278
rect 6300 800 6356 3276
rect 6524 3266 6580 3276
rect 8988 3330 9380 3332
rect 8988 3278 9326 3330
rect 9378 3278 9380 3330
rect 8988 3276 9380 3278
rect 8988 800 9044 3276
rect 9324 3266 9380 3276
rect 11676 3330 11956 3332
rect 11676 3278 11902 3330
rect 11954 3278 11956 3330
rect 11676 3276 11956 3278
rect 11676 800 11732 3276
rect 11900 3266 11956 3276
rect 14364 3330 14644 3332
rect 14364 3278 14590 3330
rect 14642 3278 14644 3330
rect 14364 3276 14644 3278
rect 14364 800 14420 3276
rect 14588 3266 14644 3276
rect 17052 3330 17332 3332
rect 17052 3278 17278 3330
rect 17330 3278 17332 3330
rect 17052 3276 17332 3278
rect 17052 800 17108 3276
rect 17276 3266 17332 3276
rect 19628 3330 20020 3332
rect 19628 3278 19966 3330
rect 20018 3278 20020 3330
rect 19628 3276 20020 3278
rect 19628 980 19684 3276
rect 19964 3266 20020 3276
rect 22428 3330 22708 3332
rect 22428 3278 22654 3330
rect 22706 3278 22708 3330
rect 22428 3276 22708 3278
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 19628 924 19796 980
rect 19740 800 19796 924
rect 22428 800 22484 3276
rect 22652 3266 22708 3276
rect 25116 3330 25396 3332
rect 25116 3278 25342 3330
rect 25394 3278 25396 3330
rect 25116 3276 25396 3278
rect 25116 800 25172 3276
rect 25340 3266 25396 3276
rect 27804 800 27860 3612
rect 28588 3668 28644 3678
rect 28588 3574 28644 3612
rect 30604 2100 30660 4062
rect 31500 3668 31556 5740
rect 33180 4564 33236 6860
rect 39228 6804 39284 6814
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 35644 4564 35700 4574
rect 32508 4562 33236 4564
rect 32508 4510 33182 4562
rect 33234 4510 33236 4562
rect 32508 4508 33236 4510
rect 32508 4338 32564 4508
rect 33180 4498 33236 4508
rect 35532 4508 35644 4564
rect 32508 4286 32510 4338
rect 32562 4286 32564 4338
rect 32508 4274 32564 4286
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 30940 3666 31556 3668
rect 30940 3614 31502 3666
rect 31554 3614 31556 3666
rect 30940 3612 31556 3614
rect 30940 3554 30996 3612
rect 31500 3602 31556 3612
rect 33180 3666 33236 3678
rect 33180 3614 33182 3666
rect 33234 3614 33236 3666
rect 30940 3502 30942 3554
rect 30994 3502 30996 3554
rect 30940 3490 30996 3502
rect 30492 2044 30660 2100
rect 30492 800 30548 2044
rect 33180 800 33236 3614
rect 35420 3556 35476 3566
rect 35532 3556 35588 4508
rect 35644 4470 35700 4508
rect 36316 3668 36372 3678
rect 39228 3668 39284 6748
rect 44492 6020 44548 6030
rect 44492 4564 44548 5964
rect 49756 5234 49812 7532
rect 50556 6300 50820 6310
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50556 6234 50820 6244
rect 49756 5182 49758 5234
rect 49810 5182 49812 5234
rect 49756 5124 49812 5182
rect 52108 5234 52164 9212
rect 52108 5182 52110 5234
rect 52162 5182 52164 5234
rect 50092 5124 50148 5134
rect 49756 5122 50148 5124
rect 49756 5070 50094 5122
rect 50146 5070 50148 5122
rect 49756 5068 50148 5070
rect 52108 5124 52164 5182
rect 55132 5236 55188 26012
rect 57820 12740 57876 12750
rect 57036 5908 57092 5918
rect 55132 5234 55524 5236
rect 55132 5182 55134 5234
rect 55186 5182 55524 5234
rect 55132 5180 55524 5182
rect 55132 5170 55188 5180
rect 52780 5124 52836 5134
rect 52108 5122 52836 5124
rect 52108 5070 52782 5122
rect 52834 5070 52836 5122
rect 52108 5068 52836 5070
rect 50092 5058 50148 5068
rect 52780 5058 52836 5068
rect 55468 5122 55524 5180
rect 55468 5070 55470 5122
rect 55522 5070 55524 5122
rect 55468 5058 55524 5070
rect 46956 4900 47012 4910
rect 46956 4564 47012 4844
rect 44044 4562 44548 4564
rect 44044 4510 44494 4562
rect 44546 4510 44548 4562
rect 44044 4508 44548 4510
rect 44044 4338 44100 4508
rect 44492 4498 44548 4508
rect 46732 4562 47012 4564
rect 46732 4510 46958 4562
rect 47010 4510 47012 4562
rect 46732 4508 47012 4510
rect 44044 4286 44046 4338
rect 44098 4286 44100 4338
rect 44044 4274 44100 4286
rect 41692 4116 41748 4126
rect 35420 3554 35588 3556
rect 35420 3502 35422 3554
rect 35474 3502 35588 3554
rect 35420 3500 35588 3502
rect 35868 3666 36372 3668
rect 35868 3614 36318 3666
rect 36370 3614 36372 3666
rect 35868 3612 36372 3614
rect 35420 3490 35476 3500
rect 35868 800 35924 3612
rect 36316 3602 36372 3612
rect 38668 3666 39284 3668
rect 38668 3614 39230 3666
rect 39282 3614 39284 3666
rect 38668 3612 39284 3614
rect 38668 3554 38724 3612
rect 39228 3602 39284 3612
rect 41244 4114 41748 4116
rect 41244 4062 41694 4114
rect 41746 4062 41748 4114
rect 41244 4060 41748 4062
rect 38668 3502 38670 3554
rect 38722 3502 38724 3554
rect 38668 3490 38724 3502
rect 38556 3444 38612 3454
rect 38556 800 38612 3388
rect 40572 3444 40628 3454
rect 40572 3350 40628 3388
rect 41244 800 41300 4060
rect 41692 4050 41748 4060
rect 42364 3668 42420 3678
rect 42364 3554 42420 3612
rect 42924 3668 42980 3678
rect 44380 3668 44436 3678
rect 42924 3574 42980 3612
rect 43932 3666 44436 3668
rect 43932 3614 44382 3666
rect 44434 3614 44436 3666
rect 43932 3612 44436 3614
rect 42364 3502 42366 3554
rect 42418 3502 42420 3554
rect 42364 3490 42420 3502
rect 43932 800 43988 3612
rect 44380 3602 44436 3612
rect 46732 3554 46788 4508
rect 46956 4498 47012 4508
rect 50428 4898 50484 4910
rect 50428 4846 50430 4898
rect 50482 4846 50484 4898
rect 49980 4228 50036 4238
rect 49756 4116 49812 4126
rect 49308 4114 49812 4116
rect 49308 4062 49758 4114
rect 49810 4062 49812 4114
rect 49308 4060 49812 4062
rect 46732 3502 46734 3554
rect 46786 3502 46788 3554
rect 46732 3490 46788 3502
rect 47628 3666 47684 3678
rect 47628 3614 47630 3666
rect 47682 3614 47684 3666
rect 46620 3444 46676 3454
rect 46620 800 46676 3388
rect 47628 3444 47684 3614
rect 47628 3378 47684 3388
rect 49308 800 49364 4060
rect 49756 4050 49812 4060
rect 49980 3554 50036 4172
rect 49980 3502 49982 3554
rect 50034 3502 50036 3554
rect 49980 3490 50036 3502
rect 50428 3556 50484 4846
rect 53116 4898 53172 4910
rect 53116 4846 53118 4898
rect 53170 4846 53172 4898
rect 50556 4732 50820 4742
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50556 4666 50820 4676
rect 51996 4452 52052 4462
rect 51996 4338 52052 4396
rect 52556 4452 52612 4462
rect 52556 4358 52612 4396
rect 51996 4286 51998 4338
rect 52050 4286 52052 4338
rect 51996 4274 52052 4286
rect 50540 4228 50596 4238
rect 50540 3666 50596 4172
rect 50540 3614 50542 3666
rect 50594 3614 50596 3666
rect 50540 3602 50596 3614
rect 52892 3666 52948 3678
rect 52892 3614 52894 3666
rect 52946 3614 52948 3666
rect 50428 3490 50484 3500
rect 51884 3556 51940 3566
rect 51884 3462 51940 3500
rect 51996 3444 52052 3454
rect 50556 3164 50820 3174
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50556 3098 50820 3108
rect 51996 800 52052 3388
rect 52892 3444 52948 3614
rect 53116 3556 53172 4846
rect 55804 4898 55860 4910
rect 55804 4846 55806 4898
rect 55858 4846 55860 4898
rect 55804 4340 55860 4846
rect 55804 4274 55860 4284
rect 57036 4228 57092 5852
rect 57820 5236 57876 12684
rect 58044 12740 58100 45836
rect 58156 45890 58212 45902
rect 58156 45838 58158 45890
rect 58210 45838 58212 45890
rect 58156 45668 58212 45838
rect 62076 45890 62132 45902
rect 62076 45838 62078 45890
rect 62130 45838 62132 45890
rect 58156 45602 58212 45612
rect 58940 45668 58996 45678
rect 58940 45574 58996 45612
rect 61292 45668 61348 45678
rect 58044 12674 58100 12684
rect 59948 14308 60004 14318
rect 59948 5236 60004 14252
rect 61292 14308 61348 45612
rect 62076 45668 62132 45838
rect 65884 45890 65940 45902
rect 65884 45838 65886 45890
rect 65938 45838 65940 45890
rect 65884 45780 65940 45838
rect 69692 45892 69748 45902
rect 69692 45890 69972 45892
rect 69692 45838 69694 45890
rect 69746 45838 69972 45890
rect 69692 45836 69972 45838
rect 69692 45826 69748 45836
rect 65884 45714 65940 45724
rect 66556 45780 66612 45790
rect 66556 45686 66612 45724
rect 62076 45602 62132 45612
rect 62748 45668 62804 45678
rect 62748 45574 62804 45612
rect 69692 45668 69748 45678
rect 65916 44716 66180 44726
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 65916 44650 66180 44660
rect 65916 43148 66180 43158
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 65916 43082 66180 43092
rect 65916 41580 66180 41590
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 65916 41514 66180 41524
rect 65916 40012 66180 40022
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 65916 39946 66180 39956
rect 65916 38444 66180 38454
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 65916 38378 66180 38388
rect 65916 36876 66180 36886
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 65916 36810 66180 36820
rect 65916 35308 66180 35318
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 65916 35242 66180 35252
rect 65916 33740 66180 33750
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 65916 33674 66180 33684
rect 65916 32172 66180 32182
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 65916 32106 66180 32116
rect 65916 30604 66180 30614
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 65916 30538 66180 30548
rect 65916 29036 66180 29046
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 65916 28970 66180 28980
rect 65916 27468 66180 27478
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 65916 27402 66180 27412
rect 65916 25900 66180 25910
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 65916 25834 66180 25844
rect 65916 24332 66180 24342
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 65916 24266 66180 24276
rect 65916 22764 66180 22774
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 65916 22698 66180 22708
rect 65916 21196 66180 21206
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 65916 21130 66180 21140
rect 65916 19628 66180 19638
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 65916 19562 66180 19572
rect 68572 19348 68628 19358
rect 65916 18060 66180 18070
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 65916 17994 66180 18004
rect 65916 16492 66180 16502
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 65916 16426 66180 16436
rect 61292 14242 61348 14252
rect 63196 15988 63252 15998
rect 57820 5234 58212 5236
rect 57820 5182 57822 5234
rect 57874 5182 58212 5234
rect 57820 5180 58212 5182
rect 57820 5170 57876 5180
rect 58156 5122 58212 5180
rect 59948 5142 60004 5180
rect 60844 5236 60900 5246
rect 58156 5070 58158 5122
rect 58210 5070 58212 5122
rect 58156 5058 58212 5070
rect 60844 5122 60900 5180
rect 63196 5236 63252 15932
rect 65916 14924 66180 14934
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 65916 14858 66180 14868
rect 65916 13356 66180 13366
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 65916 13290 66180 13300
rect 65916 11788 66180 11798
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 65916 11722 66180 11732
rect 65436 11284 65492 11294
rect 65436 5908 65492 11228
rect 65916 10220 66180 10230
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 65916 10154 66180 10164
rect 65916 8652 66180 8662
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 65916 8586 66180 8596
rect 65916 7084 66180 7094
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 65916 7018 66180 7028
rect 65436 5852 65828 5908
rect 65772 5236 65828 5852
rect 65916 5516 66180 5526
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 65916 5450 66180 5460
rect 65884 5236 65940 5246
rect 68572 5236 68628 19292
rect 69692 15988 69748 45612
rect 69916 45668 69972 45836
rect 73500 45890 73556 45902
rect 73500 45838 73502 45890
rect 73554 45838 73556 45890
rect 69916 45602 69972 45612
rect 70364 45668 70420 45678
rect 70364 45574 70420 45612
rect 73276 45668 73332 45678
rect 73276 17668 73332 45612
rect 73500 45668 73556 45838
rect 73500 45602 73556 45612
rect 74172 45668 74228 45678
rect 74172 45574 74228 45612
rect 75516 44996 75572 49200
rect 79548 46004 79604 49200
rect 83580 46004 83636 49200
rect 87612 46004 87668 49200
rect 91644 46004 91700 49200
rect 95676 46004 95732 49200
rect 99708 47012 99764 49200
rect 99708 46956 100212 47012
rect 96636 46284 96900 46294
rect 96692 46228 96740 46284
rect 96796 46228 96844 46284
rect 96636 46218 96900 46228
rect 79548 46002 79828 46004
rect 79548 45950 79550 46002
rect 79602 45950 79828 46002
rect 79548 45948 79828 45950
rect 79548 45938 79604 45948
rect 79772 45890 79828 45948
rect 83580 46002 83860 46004
rect 83580 45950 83582 46002
rect 83634 45950 83860 46002
rect 83580 45948 83860 45950
rect 83580 45938 83636 45948
rect 79772 45838 79774 45890
rect 79826 45838 79828 45890
rect 79772 45826 79828 45838
rect 83804 45890 83860 45948
rect 87612 46002 87892 46004
rect 87612 45950 87614 46002
rect 87666 45950 87892 46002
rect 87612 45948 87892 45950
rect 87612 45938 87668 45948
rect 83804 45838 83806 45890
rect 83858 45838 83860 45890
rect 83804 45826 83860 45838
rect 87836 45890 87892 45948
rect 91644 46002 91924 46004
rect 91644 45950 91646 46002
rect 91698 45950 91924 46002
rect 91644 45948 91924 45950
rect 91644 45938 91700 45948
rect 87836 45838 87838 45890
rect 87890 45838 87892 45890
rect 87836 45826 87892 45838
rect 91868 45890 91924 45948
rect 95676 46002 95956 46004
rect 95676 45950 95678 46002
rect 95730 45950 95956 46002
rect 95676 45948 95956 45950
rect 95676 45938 95732 45948
rect 91868 45838 91870 45890
rect 91922 45838 91924 45890
rect 91868 45826 91924 45838
rect 95900 45890 95956 45948
rect 95900 45838 95902 45890
rect 95954 45838 95956 45890
rect 95900 45826 95956 45838
rect 100156 46002 100212 46956
rect 100156 45950 100158 46002
rect 100210 45950 100212 46002
rect 100156 45892 100212 45950
rect 103740 46004 103796 49200
rect 103964 46004 104020 46014
rect 103740 46002 104020 46004
rect 103740 45950 103966 46002
rect 104018 45950 104020 46002
rect 103740 45948 104020 45950
rect 100156 45826 100212 45836
rect 100828 45892 100884 45902
rect 100828 45798 100884 45836
rect 103964 45892 104020 45948
rect 107772 46004 107828 49200
rect 111692 46004 111748 46014
rect 111804 46004 111860 49200
rect 115836 46900 115892 49200
rect 115500 46844 116116 46900
rect 107772 46002 108388 46004
rect 107772 45950 107774 46002
rect 107826 45950 108388 46002
rect 107772 45948 108388 45950
rect 107772 45938 107828 45948
rect 103964 45826 104020 45836
rect 104636 45892 104692 45902
rect 104636 45798 104692 45836
rect 108332 45890 108388 45948
rect 111692 46002 112196 46004
rect 111692 45950 111694 46002
rect 111746 45950 112196 46002
rect 111692 45948 112196 45950
rect 111692 45938 111748 45948
rect 108332 45838 108334 45890
rect 108386 45838 108388 45890
rect 108332 45826 108388 45838
rect 112140 45890 112196 45948
rect 115500 46002 115556 46844
rect 115500 45950 115502 46002
rect 115554 45950 115556 46002
rect 115500 45938 115556 45950
rect 112140 45838 112142 45890
rect 112194 45838 112196 45890
rect 112140 45826 112196 45838
rect 116060 45890 116116 46844
rect 119308 46004 119364 46014
rect 119868 46004 119924 49200
rect 119308 46002 119924 46004
rect 119308 45950 119310 46002
rect 119362 45950 119924 46002
rect 119308 45948 119924 45950
rect 119308 45938 119364 45948
rect 116060 45838 116062 45890
rect 116114 45838 116116 45890
rect 116060 45826 116116 45838
rect 119868 45892 119924 45948
rect 123900 46004 123956 49200
rect 127356 46284 127620 46294
rect 127412 46228 127460 46284
rect 127516 46228 127564 46284
rect 127356 46218 127620 46228
rect 127932 46004 127988 49200
rect 131964 46004 132020 49200
rect 135996 46004 136052 49200
rect 140028 46004 140084 49200
rect 144060 46004 144116 49200
rect 148092 46116 148148 49200
rect 148092 46050 148148 46060
rect 150444 46116 150500 46126
rect 150444 46022 150500 46060
rect 150332 46004 150388 46014
rect 123900 46002 124180 46004
rect 123900 45950 123902 46002
rect 123954 45950 124180 46002
rect 123900 45948 124180 45950
rect 123900 45938 123956 45948
rect 120092 45892 120148 45902
rect 119868 45890 120148 45892
rect 119868 45838 120094 45890
rect 120146 45838 120148 45890
rect 119868 45836 120148 45838
rect 120092 45826 120148 45836
rect 124124 45890 124180 45948
rect 127932 46002 128212 46004
rect 127932 45950 127934 46002
rect 127986 45950 128212 46002
rect 127932 45948 128212 45950
rect 127932 45938 127988 45948
rect 124124 45838 124126 45890
rect 124178 45838 124180 45890
rect 124124 45826 124180 45838
rect 128156 45890 128212 45948
rect 131964 46002 132244 46004
rect 131964 45950 131966 46002
rect 132018 45950 132244 46002
rect 131964 45948 132244 45950
rect 131964 45938 132020 45948
rect 128156 45838 128158 45890
rect 128210 45838 128212 45890
rect 128156 45826 128212 45838
rect 132188 45890 132244 45948
rect 135996 46002 136500 46004
rect 135996 45950 135998 46002
rect 136050 45950 136500 46002
rect 135996 45948 136500 45950
rect 135996 45938 136052 45948
rect 132188 45838 132190 45890
rect 132242 45838 132244 45890
rect 132188 45826 132244 45838
rect 136444 45890 136500 45948
rect 140028 46002 140532 46004
rect 140028 45950 140030 46002
rect 140082 45950 140532 46002
rect 140028 45948 140532 45950
rect 140028 45938 140084 45948
rect 136444 45838 136446 45890
rect 136498 45838 136500 45890
rect 136444 45826 136500 45838
rect 140476 45890 140532 45948
rect 144060 46002 144564 46004
rect 144060 45950 144062 46002
rect 144114 45950 144564 46002
rect 144060 45948 144564 45950
rect 144060 45938 144116 45948
rect 140476 45838 140478 45890
rect 140530 45838 140532 45890
rect 140476 45826 140532 45838
rect 144508 45890 144564 45948
rect 144508 45838 144510 45890
rect 144562 45838 144564 45890
rect 144508 45826 144564 45838
rect 130172 45780 130228 45790
rect 76412 45668 76468 45678
rect 75964 44996 76020 45006
rect 75516 44994 76020 44996
rect 75516 44942 75966 44994
rect 76018 44942 76020 44994
rect 75516 44940 76020 44942
rect 75964 44930 76020 44940
rect 76412 19348 76468 45612
rect 80108 45666 80164 45678
rect 80108 45614 80110 45666
rect 80162 45614 80164 45666
rect 78316 45108 78372 45118
rect 78876 45108 78932 45118
rect 78316 45106 78932 45108
rect 78316 45054 78318 45106
rect 78370 45054 78878 45106
rect 78930 45054 78932 45106
rect 78316 45052 78932 45054
rect 78316 31948 78372 45052
rect 78876 45042 78932 45052
rect 80108 43652 80164 45614
rect 84140 45666 84196 45678
rect 84140 45614 84142 45666
rect 84194 45614 84196 45666
rect 81276 45500 81540 45510
rect 81332 45444 81380 45500
rect 81436 45444 81484 45500
rect 81276 45434 81540 45444
rect 81276 43932 81540 43942
rect 81332 43876 81380 43932
rect 81436 43876 81484 43932
rect 81276 43866 81540 43876
rect 80108 43586 80164 43596
rect 81276 42364 81540 42374
rect 81332 42308 81380 42364
rect 81436 42308 81484 42364
rect 81276 42298 81540 42308
rect 81276 40796 81540 40806
rect 81332 40740 81380 40796
rect 81436 40740 81484 40796
rect 81276 40730 81540 40740
rect 81276 39228 81540 39238
rect 81332 39172 81380 39228
rect 81436 39172 81484 39228
rect 81276 39162 81540 39172
rect 81276 37660 81540 37670
rect 81332 37604 81380 37660
rect 81436 37604 81484 37660
rect 81276 37594 81540 37604
rect 81276 36092 81540 36102
rect 81332 36036 81380 36092
rect 81436 36036 81484 36092
rect 81276 36026 81540 36036
rect 84140 34692 84196 45614
rect 88172 45666 88228 45678
rect 88172 45614 88174 45666
rect 88226 45614 88228 45666
rect 88172 39508 88228 45614
rect 92204 45666 92260 45678
rect 92204 45614 92206 45666
rect 92258 45614 92260 45666
rect 92204 41188 92260 45614
rect 96236 45666 96292 45678
rect 96236 45614 96238 45666
rect 96290 45614 96292 45666
rect 96236 43708 96292 45614
rect 101052 45666 101108 45678
rect 101052 45614 101054 45666
rect 101106 45614 101108 45666
rect 96636 44716 96900 44726
rect 96692 44660 96740 44716
rect 96796 44660 96844 44716
rect 96636 44650 96900 44660
rect 101052 43708 101108 45614
rect 104860 45666 104916 45678
rect 104860 45614 104862 45666
rect 104914 45614 104916 45666
rect 104860 43708 104916 45614
rect 108668 45666 108724 45678
rect 108668 45614 108670 45666
rect 108722 45614 108724 45666
rect 96236 43652 97188 43708
rect 101052 43652 101780 43708
rect 104860 43652 105476 43708
rect 96636 43148 96900 43158
rect 96692 43092 96740 43148
rect 96796 43092 96844 43148
rect 96636 43082 96900 43092
rect 96636 41580 96900 41590
rect 96692 41524 96740 41580
rect 96796 41524 96844 41580
rect 96636 41514 96900 41524
rect 92204 41122 92260 41132
rect 96636 40012 96900 40022
rect 96692 39956 96740 40012
rect 96796 39956 96844 40012
rect 96636 39946 96900 39956
rect 88172 39442 88228 39452
rect 96636 38444 96900 38454
rect 96692 38388 96740 38444
rect 96796 38388 96844 38444
rect 96636 38378 96900 38388
rect 96636 36876 96900 36886
rect 96692 36820 96740 36876
rect 96796 36820 96844 36876
rect 96636 36810 96900 36820
rect 96636 35308 96900 35318
rect 96692 35252 96740 35308
rect 96796 35252 96844 35308
rect 96636 35242 96900 35252
rect 84140 34626 84196 34636
rect 81276 34524 81540 34534
rect 81332 34468 81380 34524
rect 81436 34468 81484 34524
rect 81276 34458 81540 34468
rect 96636 33740 96900 33750
rect 96692 33684 96740 33740
rect 96796 33684 96844 33740
rect 96636 33674 96900 33684
rect 81276 32956 81540 32966
rect 81332 32900 81380 32956
rect 81436 32900 81484 32956
rect 81276 32890 81540 32900
rect 96636 32172 96900 32182
rect 96692 32116 96740 32172
rect 96796 32116 96844 32172
rect 96636 32106 96900 32116
rect 76412 19282 76468 19292
rect 77868 31892 78372 31948
rect 73276 17602 73332 17612
rect 69692 15922 69748 15932
rect 77868 11284 77924 31892
rect 81276 31388 81540 31398
rect 81332 31332 81380 31388
rect 81436 31332 81484 31388
rect 81276 31322 81540 31332
rect 96636 30604 96900 30614
rect 96692 30548 96740 30604
rect 96796 30548 96844 30604
rect 96636 30538 96900 30548
rect 96236 30212 96292 30222
rect 96236 30118 96292 30156
rect 96684 30212 96740 30222
rect 96684 30118 96740 30156
rect 93772 30100 93828 30110
rect 81276 29820 81540 29830
rect 81332 29764 81380 29820
rect 81436 29764 81484 29820
rect 81276 29754 81540 29764
rect 81276 28252 81540 28262
rect 81332 28196 81380 28252
rect 81436 28196 81484 28252
rect 81276 28186 81540 28196
rect 81276 26684 81540 26694
rect 81332 26628 81380 26684
rect 81436 26628 81484 26684
rect 81276 26618 81540 26628
rect 81276 25116 81540 25126
rect 81332 25060 81380 25116
rect 81436 25060 81484 25116
rect 81276 25050 81540 25060
rect 81276 23548 81540 23558
rect 81332 23492 81380 23548
rect 81436 23492 81484 23548
rect 81276 23482 81540 23492
rect 81276 21980 81540 21990
rect 81332 21924 81380 21980
rect 81436 21924 81484 21980
rect 81276 21914 81540 21924
rect 81276 20412 81540 20422
rect 81332 20356 81380 20412
rect 81436 20356 81484 20412
rect 81276 20346 81540 20356
rect 81276 18844 81540 18854
rect 81332 18788 81380 18844
rect 81436 18788 81484 18844
rect 81276 18778 81540 18788
rect 81276 17276 81540 17286
rect 81332 17220 81380 17276
rect 81436 17220 81484 17276
rect 81276 17210 81540 17220
rect 81276 15708 81540 15718
rect 81332 15652 81380 15708
rect 81436 15652 81484 15708
rect 81276 15642 81540 15652
rect 81276 14140 81540 14150
rect 81332 14084 81380 14140
rect 81436 14084 81484 14140
rect 81276 14074 81540 14084
rect 81276 12572 81540 12582
rect 81332 12516 81380 12572
rect 81436 12516 81484 12572
rect 81276 12506 81540 12516
rect 77868 11218 77924 11228
rect 81276 11004 81540 11014
rect 81332 10948 81380 11004
rect 81436 10948 81484 11004
rect 81276 10938 81540 10948
rect 81276 9436 81540 9446
rect 81332 9380 81380 9436
rect 81436 9380 81484 9436
rect 81276 9370 81540 9380
rect 88060 8484 88116 8494
rect 81276 7868 81540 7878
rect 81332 7812 81380 7868
rect 81436 7812 81484 7868
rect 81276 7802 81540 7812
rect 73052 6468 73108 6478
rect 63196 5234 63588 5236
rect 63196 5182 63198 5234
rect 63250 5182 63588 5234
rect 63196 5180 63588 5182
rect 65772 5234 66276 5236
rect 65772 5182 65886 5234
rect 65938 5182 66276 5234
rect 65772 5180 66276 5182
rect 63196 5170 63252 5180
rect 60844 5070 60846 5122
rect 60898 5070 60900 5122
rect 60844 5058 60900 5070
rect 63532 5122 63588 5180
rect 65884 5170 65940 5180
rect 63532 5070 63534 5122
rect 63586 5070 63588 5122
rect 63532 5058 63588 5070
rect 66220 5122 66276 5180
rect 68572 5234 68964 5236
rect 68572 5182 68574 5234
rect 68626 5182 68964 5234
rect 68572 5180 68964 5182
rect 68572 5170 68628 5180
rect 66220 5070 66222 5122
rect 66274 5070 66276 5122
rect 66220 5058 66276 5070
rect 68908 5122 68964 5180
rect 68908 5070 68910 5122
rect 68962 5070 68964 5122
rect 68908 5058 68964 5070
rect 58492 4898 58548 4910
rect 58492 4846 58494 4898
rect 58546 4846 58548 4898
rect 57596 4340 57652 4350
rect 57596 4246 57652 4284
rect 57036 4162 57092 4172
rect 57372 4116 57428 4126
rect 56028 3668 56084 3678
rect 56028 3574 56084 3612
rect 53116 3490 53172 3500
rect 55020 3556 55076 3566
rect 55020 3462 55076 3500
rect 52892 3378 52948 3388
rect 54684 3444 54740 3454
rect 54684 800 54740 3388
rect 57372 800 57428 4060
rect 58492 3556 58548 4846
rect 61180 4898 61236 4910
rect 61180 4846 61182 4898
rect 61234 4846 61236 4898
rect 58604 4116 58660 4126
rect 58604 4022 58660 4060
rect 60508 3668 60564 3678
rect 60060 3666 60564 3668
rect 60060 3614 60510 3666
rect 60562 3614 60564 3666
rect 60060 3612 60564 3614
rect 58492 3490 58548 3500
rect 59500 3556 59556 3566
rect 59500 3462 59556 3500
rect 60060 800 60116 3612
rect 60508 3602 60564 3612
rect 61180 3556 61236 4846
rect 63868 4898 63924 4910
rect 63868 4846 63870 4898
rect 63922 4846 63924 4898
rect 61180 3490 61236 3500
rect 62748 3668 62804 3678
rect 62748 800 62804 3612
rect 62972 3556 63028 3566
rect 62972 3462 63028 3500
rect 63868 3556 63924 4846
rect 66556 4898 66612 4910
rect 66556 4846 66558 4898
rect 66610 4846 66612 4898
rect 66556 4340 66612 4846
rect 69244 4898 69300 4910
rect 69244 4846 69246 4898
rect 69298 4846 69300 4898
rect 66556 4274 66612 4284
rect 68348 4340 68404 4350
rect 68348 4246 68404 4284
rect 68124 4116 68180 4126
rect 65916 3948 66180 3958
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 65916 3882 66180 3892
rect 63980 3668 64036 3678
rect 63980 3574 64036 3612
rect 67452 3668 67508 3678
rect 67452 3574 67508 3612
rect 63868 3490 63924 3500
rect 66444 3556 66500 3566
rect 66444 3462 66500 3500
rect 65436 3444 65492 3454
rect 65436 800 65492 3388
rect 68124 800 68180 4060
rect 69244 3556 69300 4846
rect 73052 4452 73108 6412
rect 81276 6300 81540 6310
rect 81332 6244 81380 6300
rect 81436 6244 81484 6300
rect 81276 6234 81540 6244
rect 84252 5684 84308 5694
rect 81276 4732 81540 4742
rect 81332 4676 81380 4732
rect 81436 4676 81484 4732
rect 81276 4666 81540 4676
rect 73052 4386 73108 4396
rect 77196 4452 77252 4462
rect 69356 4116 69412 4126
rect 76636 4116 76692 4126
rect 69356 4022 69412 4060
rect 76188 4114 76692 4116
rect 76188 4062 76638 4114
rect 76690 4062 76692 4114
rect 76188 4060 76692 4062
rect 73500 3668 73556 3678
rect 69244 3490 69300 3500
rect 70924 3556 70980 3566
rect 70924 3462 70980 3500
rect 70812 3444 70868 3454
rect 70812 800 70868 3388
rect 71932 3444 71988 3454
rect 71932 3330 71988 3388
rect 71932 3278 71934 3330
rect 71986 3278 71988 3330
rect 71932 3266 71988 3278
rect 73500 800 73556 3612
rect 74284 3668 74340 3678
rect 74284 3574 74340 3612
rect 76188 800 76244 4060
rect 76636 4050 76692 4060
rect 76524 3668 76580 3678
rect 76524 3554 76580 3612
rect 77196 3668 77252 4396
rect 78876 4340 78932 4350
rect 78876 4246 78932 4284
rect 79548 4340 79604 4350
rect 79548 4246 79604 4284
rect 80556 4340 80612 4350
rect 81340 4340 81396 4350
rect 77196 3574 77252 3612
rect 78876 3666 78932 3678
rect 78876 3614 78878 3666
rect 78930 3614 78932 3666
rect 76524 3502 76526 3554
rect 76578 3502 76580 3554
rect 76524 3490 76580 3502
rect 78876 800 78932 3614
rect 80556 2324 80612 4284
rect 81116 4284 81340 4340
rect 81116 3554 81172 4284
rect 81340 4246 81396 4284
rect 84252 4340 84308 5628
rect 88060 4562 88116 8428
rect 92764 5796 92820 5806
rect 89068 5348 89124 5358
rect 88956 4564 89012 4574
rect 89068 4564 89124 5292
rect 92764 5234 92820 5740
rect 93772 5236 93828 30044
rect 95452 30100 95508 30110
rect 95452 30006 95508 30044
rect 97132 30100 97188 43652
rect 97132 30006 97188 30044
rect 101276 30212 101332 30222
rect 101276 29652 101332 30156
rect 100828 29650 101332 29652
rect 100828 29598 101278 29650
rect 101330 29598 101332 29650
rect 100828 29596 101332 29598
rect 100828 29426 100884 29596
rect 101276 29586 101332 29596
rect 101612 30100 101668 30110
rect 100828 29374 100830 29426
rect 100882 29374 100884 29426
rect 100828 29362 100884 29374
rect 97916 29316 97972 29326
rect 96636 29036 96900 29046
rect 96692 28980 96740 29036
rect 96796 28980 96844 29036
rect 96636 28970 96900 28980
rect 96636 27468 96900 27478
rect 96692 27412 96740 27468
rect 96796 27412 96844 27468
rect 96636 27402 96900 27412
rect 96636 25900 96900 25910
rect 96692 25844 96740 25900
rect 96796 25844 96844 25900
rect 96636 25834 96900 25844
rect 96636 24332 96900 24342
rect 96692 24276 96740 24332
rect 96796 24276 96844 24332
rect 96636 24266 96900 24276
rect 96636 22764 96900 22774
rect 96692 22708 96740 22764
rect 96796 22708 96844 22764
rect 96636 22698 96900 22708
rect 96636 21196 96900 21206
rect 96692 21140 96740 21196
rect 96796 21140 96844 21196
rect 96636 21130 96900 21140
rect 96636 19628 96900 19638
rect 96692 19572 96740 19628
rect 96796 19572 96844 19628
rect 96636 19562 96900 19572
rect 96636 18060 96900 18070
rect 96692 18004 96740 18060
rect 96796 18004 96844 18060
rect 96636 17994 96900 18004
rect 96636 16492 96900 16502
rect 96692 16436 96740 16492
rect 96796 16436 96844 16492
rect 96636 16426 96900 16436
rect 96636 14924 96900 14934
rect 96692 14868 96740 14924
rect 96796 14868 96844 14924
rect 96636 14858 96900 14868
rect 96636 13356 96900 13366
rect 96692 13300 96740 13356
rect 96796 13300 96844 13356
rect 96636 13290 96900 13300
rect 96636 11788 96900 11798
rect 96692 11732 96740 11788
rect 96796 11732 96844 11788
rect 96636 11722 96900 11732
rect 96636 10220 96900 10230
rect 96692 10164 96740 10220
rect 96796 10164 96844 10220
rect 96636 10154 96900 10164
rect 96636 8652 96900 8662
rect 96692 8596 96740 8652
rect 96796 8596 96844 8652
rect 96636 8586 96900 8596
rect 96636 7084 96900 7094
rect 96692 7028 96740 7084
rect 96796 7028 96844 7084
rect 96636 7018 96900 7028
rect 97468 6916 97524 6926
rect 96636 5516 96900 5526
rect 96692 5460 96740 5516
rect 96796 5460 96844 5516
rect 96636 5450 96900 5460
rect 92764 5182 92766 5234
rect 92818 5182 92820 5234
rect 92764 5170 92820 5182
rect 93324 5234 93828 5236
rect 93324 5182 93774 5234
rect 93826 5182 93828 5234
rect 93324 5180 93828 5182
rect 93324 5122 93380 5180
rect 93772 5170 93828 5180
rect 93996 5236 94052 5246
rect 93324 5070 93326 5122
rect 93378 5070 93380 5122
rect 93324 5058 93380 5070
rect 88060 4510 88062 4562
rect 88114 4510 88116 4562
rect 84252 4274 84308 4284
rect 87052 4340 87108 4350
rect 87052 4246 87108 4284
rect 88060 4340 88116 4510
rect 88060 4274 88116 4284
rect 88732 4562 89124 4564
rect 88732 4510 88958 4562
rect 89010 4510 89124 4562
rect 88732 4508 89124 4510
rect 84700 4116 84756 4126
rect 84252 4114 84756 4116
rect 84252 4062 84702 4114
rect 84754 4062 84756 4114
rect 84252 4060 84756 4062
rect 82012 3668 82068 3678
rect 81116 3502 81118 3554
rect 81170 3502 81172 3554
rect 81116 3490 81172 3502
rect 81788 3666 82068 3668
rect 81788 3614 82014 3666
rect 82066 3614 82068 3666
rect 81788 3612 82068 3614
rect 81276 3164 81540 3174
rect 81332 3108 81380 3164
rect 81436 3108 81484 3164
rect 81276 3098 81540 3108
rect 80556 2258 80612 2268
rect 81788 980 81844 3612
rect 82012 3602 82068 3612
rect 81564 924 81844 980
rect 81564 800 81620 924
rect 84252 800 84308 4060
rect 84700 4050 84756 4060
rect 84364 3554 84420 3566
rect 84364 3502 84366 3554
rect 84418 3502 84420 3554
rect 84364 3444 84420 3502
rect 88732 3554 88788 4508
rect 88956 4498 89012 4508
rect 93436 4340 93492 4350
rect 88732 3502 88734 3554
rect 88786 3502 88788 3554
rect 88732 3490 88788 3502
rect 90188 3780 90244 3790
rect 84364 3378 84420 3388
rect 84924 3444 84980 3454
rect 84924 3350 84980 3388
rect 86940 3442 86996 3454
rect 86940 3390 86942 3442
rect 86994 3390 86996 3442
rect 86940 800 86996 3390
rect 87388 3444 87444 3454
rect 87388 2548 87444 3388
rect 87388 2482 87444 2492
rect 89628 3444 89684 3454
rect 89852 3444 89908 3454
rect 89628 3442 89908 3444
rect 89628 3390 89630 3442
rect 89682 3390 89854 3442
rect 89906 3390 89908 3442
rect 89628 3388 89908 3390
rect 89628 800 89684 3388
rect 89852 3378 89908 3388
rect 90188 3442 90244 3724
rect 92652 3444 92708 3454
rect 93100 3444 93156 3454
rect 90188 3390 90190 3442
rect 90242 3390 90244 3442
rect 90188 3378 90244 3390
rect 92316 3442 93156 3444
rect 92316 3390 92654 3442
rect 92706 3390 93102 3442
rect 93154 3390 93156 3442
rect 92316 3388 93156 3390
rect 92316 800 92372 3388
rect 92652 3378 92708 3388
rect 93100 3378 93156 3388
rect 93436 3442 93492 4284
rect 93996 3668 94052 5180
rect 97468 5234 97524 6860
rect 97468 5182 97470 5234
rect 97522 5182 97524 5234
rect 97468 5170 97524 5182
rect 97916 5236 97972 29260
rect 100044 29316 100100 29326
rect 100044 29222 100100 29260
rect 98588 6132 98644 6142
rect 98476 6076 98588 6132
rect 98364 5236 98420 5246
rect 97916 5234 98420 5236
rect 97916 5182 98366 5234
rect 98418 5182 98420 5234
rect 97916 5180 98420 5182
rect 97916 5122 97972 5180
rect 98364 5170 98420 5180
rect 97916 5070 97918 5122
rect 97970 5070 97972 5122
rect 97916 5058 97972 5070
rect 98476 4676 98532 6076
rect 98588 6066 98644 6076
rect 101612 5236 101668 30044
rect 101724 29316 101780 43652
rect 104412 30212 104468 30222
rect 104412 30118 104468 30156
rect 104972 30212 105028 30222
rect 104972 30118 105028 30156
rect 103740 30100 103796 30110
rect 103740 30006 103796 30044
rect 105420 30100 105476 43652
rect 108668 31948 108724 45614
rect 112476 45666 112532 45678
rect 112476 45614 112478 45666
rect 112530 45614 112532 45666
rect 111996 45500 112260 45510
rect 112052 45444 112100 45500
rect 112156 45444 112204 45500
rect 111996 45434 112260 45444
rect 111996 43932 112260 43942
rect 112052 43876 112100 43932
rect 112156 43876 112204 43932
rect 111996 43866 112260 43876
rect 111996 42364 112260 42374
rect 112052 42308 112100 42364
rect 112156 42308 112204 42364
rect 111996 42298 112260 42308
rect 111996 40796 112260 40806
rect 112052 40740 112100 40796
rect 112156 40740 112204 40796
rect 111996 40730 112260 40740
rect 111996 39228 112260 39238
rect 112052 39172 112100 39228
rect 112156 39172 112204 39228
rect 111996 39162 112260 39172
rect 111996 37660 112260 37670
rect 112052 37604 112100 37660
rect 112156 37604 112204 37660
rect 111996 37594 112260 37604
rect 111996 36092 112260 36102
rect 112052 36036 112100 36092
rect 112156 36036 112204 36092
rect 111996 36026 112260 36036
rect 111996 34524 112260 34534
rect 112052 34468 112100 34524
rect 112156 34468 112204 34524
rect 111996 34458 112260 34468
rect 111996 32956 112260 32966
rect 112052 32900 112100 32956
rect 112156 32900 112204 32956
rect 111996 32890 112260 32900
rect 112476 31948 112532 45614
rect 116396 45666 116452 45678
rect 116396 45614 116398 45666
rect 116450 45614 116452 45666
rect 108220 31892 108724 31948
rect 111692 31892 112532 31948
rect 112588 32450 112644 32462
rect 112588 32398 112590 32450
rect 112642 32398 112644 32450
rect 105420 30006 105476 30044
rect 106540 30884 106596 30894
rect 101724 29222 101780 29260
rect 105532 6804 105588 6814
rect 102060 5236 102116 5246
rect 101612 5234 102116 5236
rect 101612 5182 102062 5234
rect 102114 5182 102116 5234
rect 101612 5180 102116 5182
rect 101612 5122 101668 5180
rect 102060 5170 102116 5180
rect 105532 5234 105588 6748
rect 106540 5236 106596 30828
rect 108220 30884 108276 31892
rect 108220 30790 108276 30828
rect 108892 30994 108948 31006
rect 108892 30942 108894 30994
rect 108946 30942 108948 30994
rect 108892 30884 108948 30942
rect 109452 30884 109508 30894
rect 108892 30882 109508 30884
rect 108892 30830 109454 30882
rect 109506 30830 109508 30882
rect 108892 30828 109508 30830
rect 108892 30324 108948 30828
rect 109452 30818 109508 30828
rect 109900 30884 109956 30894
rect 109900 30790 109956 30828
rect 108892 30258 108948 30268
rect 110796 30100 110852 30110
rect 110348 9044 110404 9054
rect 106764 6580 106820 6590
rect 105532 5182 105534 5234
rect 105586 5182 105588 5234
rect 105532 5170 105588 5182
rect 106092 5234 106596 5236
rect 106092 5182 106542 5234
rect 106594 5182 106596 5234
rect 106092 5180 106596 5182
rect 101612 5070 101614 5122
rect 101666 5070 101668 5122
rect 101612 5058 101668 5070
rect 106092 5122 106148 5180
rect 106540 5170 106596 5180
rect 106652 6524 106764 6580
rect 106092 5070 106094 5122
rect 106146 5070 106148 5122
rect 106092 5058 106148 5070
rect 98252 4620 98532 4676
rect 101052 5010 101108 5022
rect 101052 4958 101054 5010
rect 101106 4958 101108 5010
rect 96636 3948 96900 3958
rect 96692 3892 96740 3948
rect 96796 3892 96844 3948
rect 96636 3882 96900 3892
rect 93996 3602 94052 3612
rect 95564 3668 95620 3678
rect 93436 3390 93438 3442
rect 93490 3390 93492 3442
rect 93436 3378 93492 3390
rect 95004 3444 95060 3454
rect 95228 3444 95284 3454
rect 95004 3442 95284 3444
rect 95004 3390 95006 3442
rect 95058 3390 95230 3442
rect 95282 3390 95284 3442
rect 95004 3388 95284 3390
rect 95004 800 95060 3388
rect 95228 3378 95284 3388
rect 95564 3442 95620 3612
rect 95564 3390 95566 3442
rect 95618 3390 95620 3442
rect 95564 3378 95620 3390
rect 97692 3444 97748 3454
rect 97916 3444 97972 3454
rect 97692 3442 97972 3444
rect 97692 3390 97694 3442
rect 97746 3390 97918 3442
rect 97970 3390 97972 3442
rect 97692 3388 97972 3390
rect 97692 800 97748 3388
rect 97916 3378 97972 3388
rect 98252 3442 98308 4620
rect 101052 4564 101108 4958
rect 101052 4498 101108 4508
rect 103628 4116 103684 4126
rect 101052 3556 101108 3566
rect 98252 3390 98254 3442
rect 98306 3390 98308 3442
rect 98252 3378 98308 3390
rect 100268 3444 100324 3454
rect 100716 3444 100772 3454
rect 100268 3442 100772 3444
rect 100268 3390 100270 3442
rect 100322 3390 100718 3442
rect 100770 3390 100772 3442
rect 100268 3388 100772 3390
rect 100268 3378 100324 3388
rect 100380 800 100436 3388
rect 100716 3378 100772 3388
rect 101052 3442 101108 3500
rect 101052 3390 101054 3442
rect 101106 3390 101108 3442
rect 101052 3378 101108 3390
rect 103068 3444 103124 3454
rect 103292 3444 103348 3454
rect 103068 3442 103348 3444
rect 103068 3390 103070 3442
rect 103122 3390 103294 3442
rect 103346 3390 103348 3442
rect 103068 3388 103348 3390
rect 103068 800 103124 3388
rect 103292 3378 103348 3388
rect 103628 3442 103684 4060
rect 103628 3390 103630 3442
rect 103682 3390 103684 3442
rect 103628 3378 103684 3390
rect 105756 3444 105812 3454
rect 105980 3444 106036 3454
rect 105756 3442 106036 3444
rect 105756 3390 105758 3442
rect 105810 3390 105982 3442
rect 106034 3390 106036 3442
rect 105756 3388 106036 3390
rect 105756 800 105812 3388
rect 105980 3378 106036 3388
rect 106316 3444 106372 3454
rect 106652 3444 106708 6524
rect 106764 6514 106820 6524
rect 109228 5236 109284 5246
rect 109900 5236 109956 5246
rect 109228 5142 109284 5180
rect 109676 5180 109900 5236
rect 109004 5124 109060 5134
rect 106316 3442 106708 3444
rect 106316 3390 106318 3442
rect 106370 3390 106708 3442
rect 106316 3388 106708 3390
rect 107884 3444 107940 3454
rect 108668 3444 108724 3454
rect 107884 3442 108724 3444
rect 107884 3390 107886 3442
rect 107938 3390 108670 3442
rect 108722 3390 108724 3442
rect 107884 3388 108724 3390
rect 106316 3378 106372 3388
rect 107884 3378 107940 3388
rect 108444 800 108500 3388
rect 108668 3378 108724 3388
rect 109004 3442 109060 5068
rect 109676 5122 109732 5180
rect 109900 5170 109956 5180
rect 110348 5234 110404 8988
rect 110348 5182 110350 5234
rect 110402 5182 110404 5234
rect 110348 5170 110404 5182
rect 110796 5236 110852 30044
rect 111692 30100 111748 31892
rect 111996 31388 112260 31398
rect 112052 31332 112100 31388
rect 112156 31332 112204 31388
rect 111996 31322 112260 31332
rect 112364 30212 112420 30222
rect 112588 30212 112644 32398
rect 116396 31948 116452 45614
rect 120428 45666 120484 45678
rect 120428 45614 120430 45666
rect 120482 45614 120484 45666
rect 118412 41188 118468 41198
rect 117180 36260 117236 36270
rect 117180 32788 117236 36204
rect 116732 32786 117236 32788
rect 116732 32734 117182 32786
rect 117234 32734 117236 32786
rect 116732 32732 117236 32734
rect 116732 32562 116788 32732
rect 117180 32722 117236 32732
rect 116732 32510 116734 32562
rect 116786 32510 116788 32562
rect 116732 32498 116788 32510
rect 116060 31892 116452 31948
rect 116060 31220 116116 31892
rect 117292 31220 117348 31230
rect 116060 31218 117348 31220
rect 116060 31166 117294 31218
rect 117346 31166 117348 31218
rect 116060 31164 117348 31166
rect 113596 30884 113652 30894
rect 113372 30324 113428 30334
rect 113596 30324 113652 30828
rect 113428 30268 113652 30324
rect 116060 30882 116116 31164
rect 117292 31154 117348 31164
rect 116060 30830 116062 30882
rect 116114 30830 116116 30882
rect 113372 30230 113428 30268
rect 112420 30156 112644 30212
rect 112364 30118 112420 30156
rect 111692 30006 111748 30044
rect 112924 30100 112980 30110
rect 112924 30006 112980 30044
rect 111996 29820 112260 29830
rect 112052 29764 112100 29820
rect 112156 29764 112204 29820
rect 111996 29754 112260 29764
rect 111996 28252 112260 28262
rect 112052 28196 112100 28252
rect 112156 28196 112204 28252
rect 111996 28186 112260 28196
rect 111996 26684 112260 26694
rect 112052 26628 112100 26684
rect 112156 26628 112204 26684
rect 111996 26618 112260 26628
rect 111996 25116 112260 25126
rect 112052 25060 112100 25116
rect 112156 25060 112204 25116
rect 111996 25050 112260 25060
rect 111996 23548 112260 23558
rect 112052 23492 112100 23548
rect 112156 23492 112204 23548
rect 111996 23482 112260 23492
rect 111996 21980 112260 21990
rect 112052 21924 112100 21980
rect 112156 21924 112204 21980
rect 111996 21914 112260 21924
rect 111996 20412 112260 20422
rect 112052 20356 112100 20412
rect 112156 20356 112204 20412
rect 111996 20346 112260 20356
rect 111996 18844 112260 18854
rect 112052 18788 112100 18844
rect 112156 18788 112204 18844
rect 111996 18778 112260 18788
rect 111996 17276 112260 17286
rect 112052 17220 112100 17276
rect 112156 17220 112204 17276
rect 111996 17210 112260 17220
rect 111996 15708 112260 15718
rect 112052 15652 112100 15708
rect 112156 15652 112204 15708
rect 111996 15642 112260 15652
rect 111996 14140 112260 14150
rect 112052 14084 112100 14140
rect 112156 14084 112204 14140
rect 111996 14074 112260 14084
rect 111996 12572 112260 12582
rect 112052 12516 112100 12572
rect 112156 12516 112204 12572
rect 111996 12506 112260 12516
rect 111996 11004 112260 11014
rect 112052 10948 112100 11004
rect 112156 10948 112204 11004
rect 111996 10938 112260 10948
rect 112588 9940 112644 9950
rect 111996 9436 112260 9446
rect 112052 9380 112100 9436
rect 112156 9380 112204 9436
rect 111996 9370 112260 9380
rect 111996 7868 112260 7878
rect 112052 7812 112100 7868
rect 112156 7812 112204 7868
rect 111996 7802 112260 7812
rect 111996 6300 112260 6310
rect 112052 6244 112100 6300
rect 112156 6244 112204 6300
rect 111996 6234 112260 6244
rect 110796 5142 110852 5180
rect 109676 5070 109678 5122
rect 109730 5070 109732 5122
rect 109676 5058 109732 5070
rect 110012 5124 110068 5134
rect 110012 5030 110068 5068
rect 111996 4732 112260 4742
rect 112052 4676 112100 4732
rect 112156 4676 112204 4732
rect 111996 4666 112260 4676
rect 109004 3390 109006 3442
rect 109058 3390 109060 3442
rect 109004 3378 109060 3390
rect 111692 3444 111748 3454
rect 112140 3444 112196 3454
rect 111692 3442 112196 3444
rect 111692 3390 111694 3442
rect 111746 3390 112142 3442
rect 112194 3390 112196 3442
rect 111692 3388 112196 3390
rect 111692 2212 111748 3388
rect 112140 3378 112196 3388
rect 112476 3444 112532 3454
rect 112588 3444 112644 9884
rect 114492 9716 114548 9726
rect 113372 6020 113428 6030
rect 113372 5234 113428 5964
rect 113372 5182 113374 5234
rect 113426 5182 113428 5234
rect 113372 5170 113428 5182
rect 113932 5236 113988 5246
rect 113932 5122 113988 5180
rect 114380 5236 114436 5246
rect 114380 5142 114436 5180
rect 113932 5070 113934 5122
rect 113986 5070 113988 5122
rect 113932 5058 113988 5070
rect 112476 3442 112644 3444
rect 112476 3390 112478 3442
rect 112530 3390 112644 3442
rect 112476 3388 112644 3390
rect 113820 3444 113876 3454
rect 114044 3444 114100 3454
rect 113820 3442 114100 3444
rect 113820 3390 113822 3442
rect 113874 3390 114046 3442
rect 114098 3390 114100 3442
rect 113820 3388 114100 3390
rect 112476 3378 112532 3388
rect 111996 3164 112260 3174
rect 112052 3108 112100 3164
rect 112156 3108 112204 3164
rect 111996 3098 112260 3108
rect 111132 2156 111748 2212
rect 111132 800 111188 2156
rect 113820 800 113876 3388
rect 114044 3378 114100 3388
rect 114380 3444 114436 3454
rect 114492 3444 114548 9660
rect 116060 5236 116116 30830
rect 116732 30994 116788 31006
rect 116732 30942 116734 30994
rect 116786 30942 116788 30994
rect 116732 30884 116788 30942
rect 116732 30818 116788 30828
rect 117628 30884 117684 30894
rect 117628 30212 117684 30828
rect 118412 30884 118468 41132
rect 119308 37266 119364 37278
rect 119308 37214 119310 37266
rect 119362 37214 119364 37266
rect 118748 37156 118804 37166
rect 118748 37062 118804 37100
rect 119308 37156 119364 37214
rect 119308 37090 119364 37100
rect 118412 30818 118468 30828
rect 117964 30212 118020 30222
rect 117628 30210 118020 30212
rect 117628 30158 117630 30210
rect 117682 30158 117966 30210
rect 118018 30158 118020 30210
rect 117628 30156 118020 30158
rect 117628 30146 117684 30156
rect 117964 30146 118020 30156
rect 118748 30098 118804 30110
rect 118748 30046 118750 30098
rect 118802 30046 118804 30098
rect 118748 29988 118804 30046
rect 118748 8428 118804 29932
rect 120428 29988 120484 45614
rect 124460 45666 124516 45678
rect 124460 45614 124462 45666
rect 124514 45614 124516 45666
rect 124460 43708 124516 45614
rect 128492 45666 128548 45678
rect 128492 45614 128494 45666
rect 128546 45614 128548 45666
rect 127356 44716 127620 44726
rect 127412 44660 127460 44716
rect 127516 44660 127564 44716
rect 127356 44650 127620 44660
rect 124460 43652 124964 43708
rect 124236 37154 124292 37166
rect 124236 37102 124238 37154
rect 124290 37102 124292 37154
rect 124236 36260 124292 37102
rect 124236 36194 124292 36204
rect 120428 29922 120484 29932
rect 121324 29988 121380 29998
rect 121324 29894 121380 29932
rect 124460 29652 124516 29662
rect 124460 29426 124516 29596
rect 124460 29374 124462 29426
rect 124514 29374 124516 29426
rect 124460 29362 124516 29374
rect 118524 8372 118804 8428
rect 121772 29316 121828 29326
rect 116060 5170 116116 5180
rect 116844 5236 116900 5246
rect 116844 3780 116900 5180
rect 117628 5234 117684 5246
rect 118524 5236 118580 8372
rect 117628 5182 117630 5234
rect 117682 5182 117684 5234
rect 117628 4900 117684 5182
rect 118076 5234 118580 5236
rect 118076 5182 118526 5234
rect 118578 5182 118580 5234
rect 118076 5180 118580 5182
rect 118076 5122 118132 5180
rect 118524 5170 118580 5180
rect 121212 5908 121268 5918
rect 121212 5234 121268 5852
rect 121212 5182 121214 5234
rect 121266 5182 121268 5234
rect 121212 5170 121268 5182
rect 121772 5236 121828 29260
rect 123676 29316 123732 29326
rect 123676 29222 123732 29260
rect 124908 29316 124964 43652
rect 127356 43148 127620 43158
rect 127412 43092 127460 43148
rect 127516 43092 127564 43148
rect 127356 43082 127620 43092
rect 127356 41580 127620 41590
rect 127412 41524 127460 41580
rect 127516 41524 127564 41580
rect 127356 41514 127620 41524
rect 127356 40012 127620 40022
rect 127412 39956 127460 40012
rect 127516 39956 127564 40012
rect 127356 39946 127620 39956
rect 127356 38444 127620 38454
rect 127412 38388 127460 38444
rect 127516 38388 127564 38444
rect 127356 38378 127620 38388
rect 127356 36876 127620 36886
rect 127412 36820 127460 36876
rect 127516 36820 127564 36876
rect 127356 36810 127620 36820
rect 127356 35308 127620 35318
rect 127412 35252 127460 35308
rect 127516 35252 127564 35308
rect 127356 35242 127620 35252
rect 127356 33740 127620 33750
rect 127412 33684 127460 33740
rect 127516 33684 127564 33740
rect 127356 33674 127620 33684
rect 127356 32172 127620 32182
rect 127412 32116 127460 32172
rect 127516 32116 127564 32172
rect 127356 32106 127620 32116
rect 128492 31948 128548 45614
rect 128268 31892 128548 31948
rect 127356 30604 127620 30614
rect 127412 30548 127460 30604
rect 127516 30548 127564 30604
rect 127356 30538 127620 30548
rect 125356 30212 125412 30222
rect 125356 29652 125412 30156
rect 125356 29558 125412 29596
rect 126140 30100 126196 30110
rect 124908 29222 124964 29260
rect 125580 6468 125636 6478
rect 125132 6020 125188 6030
rect 122220 5236 122276 5246
rect 121772 5234 122276 5236
rect 121772 5182 122222 5234
rect 122274 5182 122276 5234
rect 121772 5180 122276 5182
rect 118076 5070 118078 5122
rect 118130 5070 118132 5122
rect 118076 5058 118132 5070
rect 121772 5122 121828 5180
rect 122220 5170 122276 5180
rect 121772 5070 121774 5122
rect 121826 5070 121828 5122
rect 121772 5058 121828 5070
rect 117628 4834 117684 4844
rect 120092 4228 120148 4238
rect 116844 3714 116900 3724
rect 117068 3780 117124 3790
rect 114380 3442 114548 3444
rect 114380 3390 114382 3442
rect 114434 3390 114548 3442
rect 114380 3388 114548 3390
rect 116508 3444 116564 3454
rect 116732 3444 116788 3454
rect 116508 3442 116788 3444
rect 116508 3390 116510 3442
rect 116562 3390 116734 3442
rect 116786 3390 116788 3442
rect 116508 3388 116788 3390
rect 114380 3378 114436 3388
rect 116508 800 116564 3388
rect 116732 3378 116788 3388
rect 117068 3442 117124 3724
rect 119308 3444 119364 3454
rect 119756 3444 119812 3454
rect 117068 3390 117070 3442
rect 117122 3390 117124 3442
rect 117068 3378 117124 3390
rect 119196 3442 119812 3444
rect 119196 3390 119310 3442
rect 119362 3390 119758 3442
rect 119810 3390 119812 3442
rect 119196 3388 119812 3390
rect 119196 800 119252 3388
rect 119308 3378 119364 3388
rect 119756 3378 119812 3388
rect 120092 3442 120148 4172
rect 120092 3390 120094 3442
rect 120146 3390 120148 3442
rect 120092 3378 120148 3390
rect 121884 3444 121940 3454
rect 122108 3444 122164 3454
rect 121884 3442 122164 3444
rect 121884 3390 121886 3442
rect 121938 3390 122110 3442
rect 122162 3390 122164 3442
rect 121884 3388 122164 3390
rect 121884 800 121940 3388
rect 122108 3378 122164 3388
rect 124572 3444 124628 3454
rect 124796 3444 124852 3454
rect 124572 3442 124852 3444
rect 124572 3390 124574 3442
rect 124626 3390 124798 3442
rect 124850 3390 124852 3442
rect 124572 3388 124852 3390
rect 122444 3330 122500 3342
rect 122444 3278 122446 3330
rect 122498 3278 122500 3330
rect 122444 2436 122500 3278
rect 122444 2370 122500 2380
rect 124572 800 124628 3388
rect 124796 3378 124852 3388
rect 125132 3442 125188 5964
rect 125580 5234 125636 6412
rect 125580 5182 125582 5234
rect 125634 5182 125636 5234
rect 125580 5170 125636 5182
rect 126140 5236 126196 30044
rect 128268 30100 128324 31892
rect 128940 30212 128996 30222
rect 128940 30118 128996 30156
rect 129948 30212 130004 30222
rect 129948 30118 130004 30156
rect 128268 30006 128324 30044
rect 129500 30100 129556 30110
rect 129500 30006 129556 30044
rect 127356 29036 127620 29046
rect 127412 28980 127460 29036
rect 127516 28980 127564 29036
rect 127356 28970 127620 28980
rect 127356 27468 127620 27478
rect 127412 27412 127460 27468
rect 127516 27412 127564 27468
rect 127356 27402 127620 27412
rect 127356 25900 127620 25910
rect 127412 25844 127460 25900
rect 127516 25844 127564 25900
rect 127356 25834 127620 25844
rect 127356 24332 127620 24342
rect 127412 24276 127460 24332
rect 127516 24276 127564 24332
rect 127356 24266 127620 24276
rect 127356 22764 127620 22774
rect 127412 22708 127460 22764
rect 127516 22708 127564 22764
rect 127356 22698 127620 22708
rect 127356 21196 127620 21206
rect 127412 21140 127460 21196
rect 127516 21140 127564 21196
rect 127356 21130 127620 21140
rect 127356 19628 127620 19638
rect 127412 19572 127460 19628
rect 127516 19572 127564 19628
rect 127356 19562 127620 19572
rect 127356 18060 127620 18070
rect 127412 18004 127460 18060
rect 127516 18004 127564 18060
rect 127356 17994 127620 18004
rect 127356 16492 127620 16502
rect 127412 16436 127460 16492
rect 127516 16436 127564 16492
rect 127356 16426 127620 16436
rect 127356 14924 127620 14934
rect 127412 14868 127460 14924
rect 127516 14868 127564 14924
rect 127356 14858 127620 14868
rect 127356 13356 127620 13366
rect 127412 13300 127460 13356
rect 127516 13300 127564 13356
rect 127356 13290 127620 13300
rect 127356 11788 127620 11798
rect 127412 11732 127460 11788
rect 127516 11732 127564 11788
rect 127356 11722 127620 11732
rect 127356 10220 127620 10230
rect 127412 10164 127460 10220
rect 127516 10164 127564 10220
rect 127356 10154 127620 10164
rect 127356 8652 127620 8662
rect 127412 8596 127460 8652
rect 127516 8596 127564 8652
rect 127356 8586 127620 8596
rect 130172 8372 130228 45724
rect 132524 45668 132580 45678
rect 136220 45668 136276 45678
rect 132524 45666 132692 45668
rect 132524 45614 132526 45666
rect 132578 45614 132692 45666
rect 132524 45612 132692 45614
rect 132524 45602 132580 45612
rect 132636 44434 132692 45612
rect 136108 45666 136276 45668
rect 136108 45614 136222 45666
rect 136274 45614 136276 45666
rect 136108 45612 136276 45614
rect 136108 45444 136164 45612
rect 136220 45602 136276 45612
rect 139916 45668 139972 45678
rect 135884 45388 136164 45444
rect 135660 45220 135716 45230
rect 135212 44994 135268 45006
rect 135212 44942 135214 44994
rect 135266 44942 135268 44994
rect 132636 44382 132638 44434
rect 132690 44382 132692 44434
rect 132636 44370 132692 44382
rect 134764 44434 134820 44446
rect 134764 44382 134766 44434
rect 134818 44382 134820 44434
rect 131964 44324 132020 44334
rect 131964 44230 132020 44268
rect 134764 42756 134820 44382
rect 135100 44324 135156 44334
rect 135212 44324 135268 44942
rect 135156 44268 135268 44324
rect 135100 43428 135156 44268
rect 135660 43708 135716 45164
rect 135884 44434 135940 45388
rect 138124 44996 138180 45006
rect 138124 44902 138180 44940
rect 138684 44996 138740 45006
rect 139692 44996 139748 45006
rect 138684 44994 138964 44996
rect 138684 44942 138686 44994
rect 138738 44942 138964 44994
rect 138684 44940 138964 44942
rect 135884 44382 135886 44434
rect 135938 44382 135940 44434
rect 135884 44370 135940 44382
rect 138012 44434 138068 44446
rect 138012 44382 138014 44434
rect 138066 44382 138068 44434
rect 138012 43708 138068 44382
rect 135660 43652 135940 43708
rect 135884 43650 135940 43652
rect 135884 43598 135886 43650
rect 135938 43598 135940 43650
rect 135884 43586 135940 43598
rect 136108 43650 136164 43662
rect 136108 43598 136110 43650
rect 136162 43598 136164 43650
rect 135772 43540 135828 43550
rect 135772 43446 135828 43484
rect 136108 43540 136164 43598
rect 137788 43652 138068 43708
rect 136108 43474 136164 43484
rect 136220 43538 136276 43550
rect 136220 43486 136222 43538
rect 136274 43486 136276 43538
rect 135100 43334 135156 43372
rect 135996 43428 136052 43438
rect 134764 42690 134820 42700
rect 133980 39508 134036 39518
rect 131068 36482 131124 36494
rect 131068 36430 131070 36482
rect 131122 36430 131124 36482
rect 130508 36260 130564 36270
rect 130508 36166 130564 36204
rect 131068 36260 131124 36430
rect 131068 36194 131124 36204
rect 132636 34692 132692 34702
rect 132636 30210 132692 34636
rect 132636 30158 132638 30210
rect 132690 30158 132692 30210
rect 132636 30100 132692 30158
rect 132860 30212 132916 30222
rect 132860 30118 132916 30156
rect 132636 30034 132692 30044
rect 133644 30100 133700 30110
rect 133644 30006 133700 30044
rect 133980 29652 134036 39452
rect 135996 36370 136052 43372
rect 136220 42532 136276 43486
rect 137228 43428 137284 43438
rect 137228 43334 137284 43372
rect 137564 43426 137620 43438
rect 137564 43374 137566 43426
rect 137618 43374 137620 43426
rect 137564 42980 137620 43374
rect 137564 42914 137620 42924
rect 137788 42978 137844 43652
rect 138684 43540 138740 44940
rect 138908 44322 138964 44940
rect 138908 44270 138910 44322
rect 138962 44270 138964 44322
rect 138908 44258 138964 44270
rect 139580 44994 139748 44996
rect 139580 44942 139694 44994
rect 139746 44942 139748 44994
rect 139580 44940 139748 44942
rect 138684 43474 138740 43484
rect 137788 42926 137790 42978
rect 137842 42926 137844 42978
rect 137788 42914 137844 42926
rect 138124 42980 138180 42990
rect 138124 42886 138180 42924
rect 137900 42756 137956 42766
rect 137900 42662 137956 42700
rect 136220 42466 136276 42476
rect 137788 42532 137844 42542
rect 137788 42438 137844 42476
rect 135996 36318 135998 36370
rect 136050 36318 136052 36370
rect 135996 35252 136052 36318
rect 136108 35252 136164 35262
rect 135996 35196 136108 35252
rect 136108 35186 136164 35196
rect 136780 35252 136836 35262
rect 136332 30884 136388 30894
rect 136332 30790 136388 30828
rect 136780 30884 136836 35196
rect 137340 30994 137396 31006
rect 137340 30942 137342 30994
rect 137394 30942 137396 30994
rect 137340 30884 137396 30942
rect 136780 30882 137396 30884
rect 136780 30830 136782 30882
rect 136834 30830 137396 30882
rect 136780 30828 137396 30830
rect 138124 30884 138180 30894
rect 135772 30324 135828 30334
rect 135772 30322 135940 30324
rect 135772 30270 135774 30322
rect 135826 30270 135940 30322
rect 135772 30268 135940 30270
rect 135772 30258 135828 30268
rect 133980 29558 134036 29596
rect 134428 30212 134484 30222
rect 134428 29652 134484 30156
rect 135772 29652 135828 29662
rect 134428 29650 135044 29652
rect 134428 29598 134430 29650
rect 134482 29598 135044 29650
rect 134428 29596 135044 29598
rect 134428 29586 134484 29596
rect 134988 29426 135044 29596
rect 135772 29538 135828 29596
rect 135772 29486 135774 29538
rect 135826 29486 135828 29538
rect 135772 29474 135828 29486
rect 134988 29374 134990 29426
rect 135042 29374 135044 29426
rect 134988 29362 135044 29374
rect 134652 17668 134708 17678
rect 132748 15988 132804 15998
rect 131068 11284 131124 11294
rect 131068 9156 131124 11228
rect 131068 9090 131124 9100
rect 130172 8306 130228 8316
rect 132748 7698 132804 15932
rect 134540 9044 134596 9054
rect 134540 8950 134596 8988
rect 132860 8372 132916 8382
rect 132860 8278 132916 8316
rect 132748 7646 132750 7698
rect 132802 7646 132804 7698
rect 132748 7634 132804 7646
rect 133084 8258 133140 8270
rect 133084 8206 133086 8258
rect 133138 8206 133140 8258
rect 132524 7588 132580 7598
rect 132524 7494 132580 7532
rect 130508 7476 130564 7486
rect 127356 7084 127620 7094
rect 127412 7028 127460 7084
rect 127516 7028 127564 7084
rect 127356 7018 127620 7028
rect 130060 6132 130116 6142
rect 127356 5516 127620 5526
rect 127412 5460 127460 5516
rect 127516 5460 127564 5516
rect 127356 5450 127620 5460
rect 126588 5236 126644 5246
rect 126140 5234 126644 5236
rect 126140 5182 126590 5234
rect 126642 5182 126644 5234
rect 126140 5180 126644 5182
rect 126140 5122 126196 5180
rect 126588 5170 126644 5180
rect 130060 5236 130116 6076
rect 130508 5346 130564 7420
rect 131740 7476 131796 7486
rect 131740 7382 131796 7420
rect 131964 7476 132020 7486
rect 131740 6916 131796 6926
rect 130508 5294 130510 5346
rect 130562 5294 130564 5346
rect 130508 5282 130564 5294
rect 131292 6692 131348 6702
rect 131292 5346 131348 6636
rect 131292 5294 131294 5346
rect 131346 5294 131348 5346
rect 131292 5282 131348 5294
rect 131740 5346 131796 6860
rect 131740 5294 131742 5346
rect 131794 5294 131796 5346
rect 131740 5282 131796 5294
rect 130396 5236 130452 5246
rect 130060 5234 130452 5236
rect 130060 5182 130062 5234
rect 130114 5182 130398 5234
rect 130450 5182 130452 5234
rect 130060 5180 130452 5182
rect 130060 5170 130116 5180
rect 130396 5170 130452 5180
rect 126140 5070 126142 5122
rect 126194 5070 126196 5122
rect 126140 5058 126196 5070
rect 131180 5122 131236 5134
rect 131180 5070 131182 5122
rect 131234 5070 131236 5122
rect 127820 4676 127876 4686
rect 127356 3948 127620 3958
rect 127412 3892 127460 3948
rect 127516 3892 127564 3948
rect 127356 3882 127620 3892
rect 125132 3390 125134 3442
rect 125186 3390 125188 3442
rect 125132 3378 125188 3390
rect 126924 3444 126980 3454
rect 127484 3444 127540 3454
rect 126924 3442 127540 3444
rect 126924 3390 126926 3442
rect 126978 3390 127486 3442
rect 127538 3390 127540 3442
rect 126924 3388 127540 3390
rect 126924 2212 126980 3388
rect 127484 3378 127540 3388
rect 127820 3442 127876 4620
rect 130508 4564 130564 4574
rect 127820 3390 127822 3442
rect 127874 3390 127876 3442
rect 127820 3378 127876 3390
rect 129948 3444 130004 3454
rect 130172 3444 130228 3454
rect 129948 3442 130228 3444
rect 129948 3390 129950 3442
rect 130002 3390 130174 3442
rect 130226 3390 130228 3442
rect 129948 3388 130228 3390
rect 126924 2156 127316 2212
rect 127260 800 127316 2156
rect 129948 800 130004 3388
rect 130172 3378 130228 3388
rect 130508 3442 130564 4508
rect 130844 4228 130900 4238
rect 131180 4228 131236 5070
rect 131628 5010 131684 5022
rect 131628 4958 131630 5010
rect 131682 4958 131684 5010
rect 130844 4226 131236 4228
rect 130844 4174 130846 4226
rect 130898 4174 131236 4226
rect 130844 4172 131236 4174
rect 131292 4228 131348 4238
rect 131628 4228 131684 4958
rect 131964 5012 132020 7420
rect 133084 6916 133140 8206
rect 134316 8260 134372 8270
rect 133084 6850 133140 6860
rect 133196 8146 133252 8158
rect 133196 8094 133198 8146
rect 133250 8094 133252 8146
rect 133196 7588 133252 8094
rect 133084 6692 133140 6702
rect 133084 6598 133140 6636
rect 132076 6580 132132 6590
rect 132076 5236 132132 6524
rect 133196 6578 133252 7532
rect 133196 6526 133198 6578
rect 133250 6526 133252 6578
rect 133196 6514 133252 6526
rect 133980 7586 134036 7598
rect 133980 7534 133982 7586
rect 134034 7534 134036 7586
rect 133756 6132 133812 6142
rect 133756 5346 133812 6076
rect 133980 5908 134036 7534
rect 134204 7474 134260 7486
rect 134204 7422 134206 7474
rect 134258 7422 134260 7474
rect 134204 6916 134260 7422
rect 134204 6850 134260 6860
rect 133980 5842 134036 5852
rect 133756 5294 133758 5346
rect 133810 5294 133812 5346
rect 133756 5282 133812 5294
rect 134204 5348 134260 5358
rect 134316 5348 134372 8204
rect 134204 5346 134372 5348
rect 134204 5294 134206 5346
rect 134258 5294 134372 5346
rect 134204 5292 134372 5294
rect 134540 7588 134596 7598
rect 134540 5346 134596 7532
rect 134652 6466 134708 17612
rect 135884 10500 135940 30268
rect 136220 30212 136276 30222
rect 136220 30118 136276 30156
rect 136780 30212 136836 30828
rect 138124 30790 138180 30828
rect 136780 30146 136836 30156
rect 137900 29314 137956 29326
rect 137900 29262 137902 29314
rect 137954 29262 137956 29314
rect 135884 10434 135940 10444
rect 136220 19348 136276 19358
rect 135324 9156 135380 9166
rect 135324 9062 135380 9100
rect 135996 9156 136052 9166
rect 135996 9062 136052 9100
rect 135548 9044 135604 9054
rect 135548 8950 135604 8988
rect 135548 8258 135604 8270
rect 135548 8206 135550 8258
rect 135602 8206 135604 8258
rect 135548 8036 135604 8206
rect 135772 8148 135828 8158
rect 135772 8054 135828 8092
rect 135548 7970 135604 7980
rect 136220 7698 136276 19292
rect 137900 11508 137956 29262
rect 139580 20188 139636 44940
rect 139692 44930 139748 44940
rect 139804 44996 139860 45006
rect 139804 44902 139860 44940
rect 139692 44436 139748 44446
rect 139916 44436 139972 45612
rect 139692 44434 139972 44436
rect 139692 44382 139694 44434
rect 139746 44382 139972 44434
rect 139692 44380 139972 44382
rect 140252 45666 140308 45678
rect 140252 45614 140254 45666
rect 140306 45614 140308 45666
rect 139692 44370 139748 44380
rect 140252 43708 140308 45614
rect 144284 45668 144340 45678
rect 144284 45574 144340 45612
rect 142716 45500 142980 45510
rect 142772 45444 142820 45500
rect 142876 45444 142924 45500
rect 142716 45434 142980 45444
rect 140588 45220 140644 45230
rect 140588 45126 140644 45164
rect 141596 45106 141652 45118
rect 141596 45054 141598 45106
rect 141650 45054 141652 45106
rect 141596 44436 141652 45054
rect 141932 44996 141988 45006
rect 141820 44436 141876 44446
rect 141596 44434 141876 44436
rect 141596 44382 141822 44434
rect 141874 44382 141876 44434
rect 141596 44380 141876 44382
rect 141820 44370 141876 44380
rect 139692 43652 140308 43708
rect 139692 43650 139748 43652
rect 139692 43598 139694 43650
rect 139746 43598 139748 43650
rect 139692 43586 139748 43598
rect 140364 43540 140420 43550
rect 140364 43446 140420 43484
rect 140252 30882 140308 30894
rect 140252 30830 140254 30882
rect 140306 30830 140308 30882
rect 139580 20132 139860 20188
rect 137900 11442 137956 11452
rect 138012 14308 138068 14318
rect 137676 10388 137732 10398
rect 137676 9042 137732 10332
rect 137676 8990 137678 9042
rect 137730 8990 137732 9042
rect 137676 8978 137732 8990
rect 136332 8148 136388 8158
rect 136332 8036 136388 8092
rect 136332 8034 136612 8036
rect 136332 7982 136334 8034
rect 136386 7982 136612 8034
rect 136332 7980 136612 7982
rect 136332 7970 136388 7980
rect 136220 7646 136222 7698
rect 136274 7646 136276 7698
rect 136220 7634 136276 7646
rect 135660 7588 135716 7598
rect 135660 7494 135716 7532
rect 135548 7476 135604 7486
rect 135548 7382 135604 7420
rect 134652 6414 134654 6466
rect 134706 6414 134708 6466
rect 134652 6402 134708 6414
rect 135212 6690 135268 6702
rect 135212 6638 135214 6690
rect 135266 6638 135268 6690
rect 134540 5294 134542 5346
rect 134594 5294 134596 5346
rect 134204 5282 134260 5292
rect 134540 5282 134596 5294
rect 135100 5908 135156 5918
rect 135100 5794 135156 5852
rect 135100 5742 135102 5794
rect 135154 5742 135156 5794
rect 132636 5236 132692 5246
rect 132076 5234 132692 5236
rect 132076 5182 132078 5234
rect 132130 5182 132638 5234
rect 132690 5182 132692 5234
rect 132076 5180 132692 5182
rect 132076 5170 132132 5180
rect 132636 5170 132692 5180
rect 133420 5236 133476 5246
rect 133476 5180 133700 5236
rect 133420 5142 133476 5180
rect 133644 5122 133700 5180
rect 133644 5070 133646 5122
rect 133698 5070 133700 5122
rect 133644 5058 133700 5070
rect 132188 5012 132244 5022
rect 131964 5010 132244 5012
rect 131964 4958 132190 5010
rect 132242 4958 132244 5010
rect 131964 4956 132244 4958
rect 132188 4946 132244 4956
rect 134092 5010 134148 5022
rect 134092 4958 134094 5010
rect 134146 4958 134148 5010
rect 131292 4226 131684 4228
rect 131292 4174 131294 4226
rect 131346 4174 131684 4226
rect 131292 4172 131684 4174
rect 132972 4340 133028 4350
rect 130844 4116 130900 4172
rect 130844 4050 130900 4060
rect 131292 3556 131348 4172
rect 132972 4116 133028 4284
rect 132972 4050 133028 4060
rect 133196 4340 133252 4350
rect 131292 3490 131348 3500
rect 130508 3390 130510 3442
rect 130562 3390 130564 3442
rect 130508 3378 130564 3390
rect 132636 3444 132692 3454
rect 132860 3444 132916 3454
rect 132636 3442 132916 3444
rect 132636 3390 132638 3442
rect 132690 3390 132862 3442
rect 132914 3390 132916 3442
rect 132636 3388 132916 3390
rect 132636 800 132692 3388
rect 132860 3378 132916 3388
rect 133196 3442 133252 4284
rect 133756 4228 133812 4238
rect 134092 4228 134148 4958
rect 133756 4226 134148 4228
rect 133756 4174 133758 4226
rect 133810 4174 134148 4226
rect 133756 4172 134148 4174
rect 133756 4116 133812 4172
rect 133756 4050 133812 4060
rect 133196 3390 133198 3442
rect 133250 3390 133252 3442
rect 133196 3378 133252 3390
rect 135100 2996 135156 5742
rect 135212 4788 135268 6638
rect 135548 6692 135604 6702
rect 135548 6132 135604 6636
rect 136332 6692 136388 6702
rect 136332 6598 136388 6636
rect 135772 6578 135828 6590
rect 135772 6526 135774 6578
rect 135826 6526 135828 6578
rect 135772 6468 135828 6526
rect 135772 6402 135828 6412
rect 135324 6130 135604 6132
rect 135324 6078 135550 6130
rect 135602 6078 135604 6130
rect 135324 6076 135604 6078
rect 135324 5122 135380 6076
rect 135548 6066 135604 6076
rect 136444 5906 136500 5918
rect 136444 5854 136446 5906
rect 136498 5854 136500 5906
rect 135772 5348 135828 5358
rect 135772 5254 135828 5292
rect 136444 5348 136500 5854
rect 136444 5282 136500 5292
rect 135324 5070 135326 5122
rect 135378 5070 135380 5122
rect 135324 5058 135380 5070
rect 135660 5010 135716 5022
rect 135660 4958 135662 5010
rect 135714 4958 135716 5010
rect 135324 4788 135380 4798
rect 135212 4732 135324 4788
rect 135324 4722 135380 4732
rect 135324 4228 135380 4238
rect 135660 4228 135716 4958
rect 135324 4226 135716 4228
rect 135324 4174 135326 4226
rect 135378 4174 135716 4226
rect 135324 4172 135716 4174
rect 135884 5012 135940 5022
rect 135324 3668 135380 4172
rect 135324 3602 135380 3612
rect 135100 2930 135156 2940
rect 135324 3444 135380 3454
rect 135548 3444 135604 3454
rect 135324 3442 135604 3444
rect 135324 3390 135326 3442
rect 135378 3390 135550 3442
rect 135602 3390 135604 3442
rect 135324 3388 135604 3390
rect 135324 800 135380 3388
rect 135548 3378 135604 3388
rect 135884 3442 135940 4956
rect 136444 4898 136500 4910
rect 136444 4846 136446 4898
rect 136498 4846 136500 4898
rect 136444 4452 136500 4846
rect 136444 4386 136500 4396
rect 135884 3390 135886 3442
rect 135938 3390 135940 3442
rect 135884 3378 135940 3390
rect 136556 2772 136612 7980
rect 137676 7588 137732 7598
rect 137676 7474 137732 7532
rect 137676 7422 137678 7474
rect 137730 7422 137732 7474
rect 137676 7410 137732 7422
rect 137228 6804 137284 6814
rect 137228 6690 137284 6748
rect 137228 6638 137230 6690
rect 137282 6638 137284 6690
rect 137228 6020 137284 6638
rect 137900 6468 137956 6478
rect 137900 6374 137956 6412
rect 138012 6130 138068 14252
rect 139132 11620 139188 11630
rect 138460 10836 138516 10846
rect 138236 10164 138292 10174
rect 138124 9156 138180 9166
rect 138124 6692 138180 9100
rect 138236 9154 138292 10108
rect 138236 9102 138238 9154
rect 138290 9102 138292 9154
rect 138236 9090 138292 9102
rect 138460 8034 138516 10780
rect 139132 10164 139188 11564
rect 138684 10052 138740 10062
rect 138684 9266 138740 9996
rect 139132 9938 139188 10108
rect 139804 10050 139860 20132
rect 140252 13524 140308 30830
rect 140252 13458 140308 13468
rect 140140 12740 140196 12750
rect 139804 9998 139806 10050
rect 139858 9998 139860 10050
rect 139804 9940 139860 9998
rect 139132 9886 139134 9938
rect 139186 9886 139188 9938
rect 139132 9874 139188 9886
rect 139580 9938 139860 9940
rect 139580 9886 139806 9938
rect 139858 9886 139860 9938
rect 139580 9884 139860 9886
rect 138684 9214 138686 9266
rect 138738 9214 138740 9266
rect 138684 9156 138740 9214
rect 139580 9266 139636 9884
rect 139804 9874 139860 9884
rect 140028 11172 140084 11182
rect 139580 9214 139582 9266
rect 139634 9214 139636 9266
rect 139580 9202 139636 9214
rect 138684 9090 138740 9100
rect 139132 9156 139188 9166
rect 139132 8930 139188 9100
rect 139132 8878 139134 8930
rect 139186 8878 139188 8930
rect 139132 8866 139188 8878
rect 139804 9156 139860 9166
rect 139468 8260 139524 8270
rect 139468 8166 139524 8204
rect 138460 7982 138462 8034
rect 138514 7982 138516 8034
rect 138236 7588 138292 7598
rect 138460 7588 138516 7982
rect 139580 8146 139636 8158
rect 139580 8094 139582 8146
rect 139634 8094 139636 8146
rect 138236 7586 138516 7588
rect 138236 7534 138238 7586
rect 138290 7534 138516 7586
rect 138236 7532 138516 7534
rect 139468 7588 139524 7598
rect 139580 7588 139636 8094
rect 139468 7586 139636 7588
rect 139468 7534 139470 7586
rect 139522 7534 139636 7586
rect 139468 7532 139636 7534
rect 138236 7522 138292 7532
rect 139132 7474 139188 7486
rect 139132 7422 139134 7474
rect 139186 7422 139188 7474
rect 138236 6692 138292 6702
rect 138124 6636 138236 6692
rect 138236 6598 138292 6636
rect 139020 6690 139076 6702
rect 139020 6638 139022 6690
rect 139074 6638 139076 6690
rect 138012 6078 138014 6130
rect 138066 6078 138068 6130
rect 138012 6066 138068 6078
rect 138908 6466 138964 6478
rect 138908 6414 138910 6466
rect 138962 6414 138964 6466
rect 136892 6018 137284 6020
rect 136892 5966 137230 6018
rect 137282 5966 137284 6018
rect 136892 5964 137284 5966
rect 136892 5122 136948 5964
rect 137228 5954 137284 5964
rect 138908 5906 138964 6414
rect 138908 5854 138910 5906
rect 138962 5854 138964 5906
rect 138908 5842 138964 5854
rect 137452 5236 137508 5246
rect 137452 5142 137508 5180
rect 136892 5070 136894 5122
rect 136946 5070 136948 5122
rect 136892 5058 136948 5070
rect 138124 5124 138180 5134
rect 138124 5030 138180 5068
rect 138908 5122 138964 5134
rect 138908 5070 138910 5122
rect 138962 5070 138964 5122
rect 137004 5010 137060 5022
rect 137004 4958 137006 5010
rect 137058 4958 137060 5010
rect 137004 4900 137060 4958
rect 137004 4834 137060 4844
rect 138012 5010 138068 5022
rect 138012 4958 138014 5010
rect 138066 4958 138068 5010
rect 138012 4900 138068 4958
rect 138908 5012 138964 5070
rect 139020 5012 139076 6638
rect 139132 6132 139188 7422
rect 139132 6066 139188 6076
rect 139244 7476 139300 7486
rect 139132 5908 139188 5918
rect 139132 5814 139188 5852
rect 139020 4956 139188 5012
rect 138908 4946 138964 4956
rect 138012 4676 138068 4844
rect 138796 4900 138852 4910
rect 138124 4676 138180 4686
rect 138012 4620 138124 4676
rect 138124 4610 138180 4620
rect 138796 4450 138852 4844
rect 138796 4398 138798 4450
rect 138850 4398 138852 4450
rect 138796 4386 138852 4398
rect 137340 4340 137396 4350
rect 137340 4246 137396 4284
rect 136556 2706 136612 2716
rect 138348 3444 138404 3454
rect 138796 3444 138852 3454
rect 138348 3442 138852 3444
rect 138348 3390 138350 3442
rect 138402 3390 138798 3442
rect 138850 3390 138852 3442
rect 138348 3388 138852 3390
rect 138348 2212 138404 3388
rect 138796 3378 138852 3388
rect 139132 3442 139188 4956
rect 139244 4562 139300 7420
rect 139468 6804 139524 7532
rect 139468 6738 139524 6748
rect 139244 4510 139246 4562
rect 139298 4510 139300 4562
rect 139244 4498 139300 4510
rect 139356 6468 139412 6478
rect 139132 3390 139134 3442
rect 139186 3390 139188 3442
rect 139132 3378 139188 3390
rect 139356 2884 139412 6412
rect 139804 6018 139860 9100
rect 140028 7698 140084 11116
rect 140140 8034 140196 12684
rect 140364 10050 140420 10062
rect 140364 9998 140366 10050
rect 140418 9998 140420 10050
rect 140364 9940 140420 9998
rect 140364 9938 140756 9940
rect 140364 9886 140366 9938
rect 140418 9886 140756 9938
rect 140364 9884 140756 9886
rect 140364 9874 140420 9884
rect 140700 9826 140756 9884
rect 140700 9774 140702 9826
rect 140754 9774 140756 9826
rect 140700 9762 140756 9774
rect 141484 9602 141540 9614
rect 141484 9550 141486 9602
rect 141538 9550 141540 9602
rect 140924 9268 140980 9278
rect 140252 9156 140308 9166
rect 140252 9062 140308 9100
rect 140924 9154 140980 9212
rect 140924 9102 140926 9154
rect 140978 9102 140980 9154
rect 140924 9090 140980 9102
rect 140140 7982 140142 8034
rect 140194 7982 140196 8034
rect 140140 7970 140196 7982
rect 140812 9042 140868 9054
rect 140812 8990 140814 9042
rect 140866 8990 140868 9042
rect 140028 7646 140030 7698
rect 140082 7646 140084 7698
rect 140028 7634 140084 7646
rect 140812 7700 140868 8990
rect 140812 7634 140868 7644
rect 140924 8258 140980 8270
rect 140924 8206 140926 8258
rect 140978 8206 140980 8258
rect 140588 7476 140644 7486
rect 140588 7382 140644 7420
rect 140364 6580 140420 6590
rect 139804 5966 139806 6018
rect 139858 5966 139860 6018
rect 139468 5796 139524 5806
rect 139468 5702 139524 5740
rect 139804 4676 139860 5966
rect 140140 6524 140364 6580
rect 140140 5906 140196 6524
rect 140140 5854 140142 5906
rect 140194 5854 140196 5906
rect 140140 5842 140196 5854
rect 140364 5010 140420 6524
rect 140700 6578 140756 6590
rect 140700 6526 140702 6578
rect 140754 6526 140756 6578
rect 140588 5796 140644 5806
rect 140588 5702 140644 5740
rect 140364 4958 140366 5010
rect 140418 4958 140420 5010
rect 140364 4900 140420 4958
rect 140364 4834 140420 4844
rect 140476 5124 140532 5134
rect 140476 5012 140532 5068
rect 140700 5012 140756 6526
rect 140476 5010 140756 5012
rect 140476 4958 140702 5010
rect 140754 4958 140756 5010
rect 140476 4956 140756 4958
rect 139804 4610 139860 4620
rect 140252 4338 140308 4350
rect 140252 4286 140254 4338
rect 140306 4286 140308 4338
rect 140252 4228 140308 4286
rect 140476 4338 140532 4956
rect 140700 4946 140756 4956
rect 140812 4900 140868 4910
rect 140924 4900 140980 8206
rect 140812 4898 140980 4900
rect 140812 4846 140814 4898
rect 140866 4846 140980 4898
rect 140812 4844 140980 4846
rect 141036 5796 141092 5806
rect 140812 4834 140868 4844
rect 140476 4286 140478 4338
rect 140530 4286 140532 4338
rect 140476 4274 140532 4286
rect 140924 4338 140980 4350
rect 140924 4286 140926 4338
rect 140978 4286 140980 4338
rect 140252 4162 140308 4172
rect 140924 3668 140980 4286
rect 140924 3602 140980 3612
rect 139356 2818 139412 2828
rect 140700 3444 140756 3454
rect 140924 3444 140980 3454
rect 140700 3442 140980 3444
rect 140700 3390 140702 3442
rect 140754 3390 140926 3442
rect 140978 3390 140980 3442
rect 140700 3388 140980 3390
rect 138012 2156 138404 2212
rect 138012 800 138068 2156
rect 140700 800 140756 3388
rect 140924 3378 140980 3388
rect 141036 2660 141092 5740
rect 141260 5794 141316 5806
rect 141260 5742 141262 5794
rect 141314 5742 141316 5794
rect 141260 5124 141316 5742
rect 141260 5058 141316 5068
rect 141484 5012 141540 9550
rect 141932 9268 141988 44940
rect 142716 43932 142980 43942
rect 142772 43876 142820 43932
rect 142876 43876 142924 43932
rect 142716 43866 142980 43876
rect 142716 42364 142980 42374
rect 142772 42308 142820 42364
rect 142876 42308 142924 42364
rect 142716 42298 142980 42308
rect 142716 40796 142980 40806
rect 142772 40740 142820 40796
rect 142876 40740 142924 40796
rect 142716 40730 142980 40740
rect 142716 39228 142980 39238
rect 142772 39172 142820 39228
rect 142876 39172 142924 39228
rect 142716 39162 142980 39172
rect 142716 37660 142980 37670
rect 142772 37604 142820 37660
rect 142876 37604 142924 37660
rect 142716 37594 142980 37604
rect 142716 36092 142980 36102
rect 142772 36036 142820 36092
rect 142876 36036 142924 36092
rect 142716 36026 142980 36036
rect 142716 34524 142980 34534
rect 142772 34468 142820 34524
rect 142876 34468 142924 34524
rect 142716 34458 142980 34468
rect 142716 32956 142980 32966
rect 142772 32900 142820 32956
rect 142876 32900 142924 32956
rect 142716 32890 142980 32900
rect 142716 31388 142980 31398
rect 142772 31332 142820 31388
rect 142876 31332 142924 31388
rect 142716 31322 142980 31332
rect 142716 29820 142980 29830
rect 142772 29764 142820 29820
rect 142876 29764 142924 29820
rect 142716 29754 142980 29764
rect 142716 28252 142980 28262
rect 142772 28196 142820 28252
rect 142876 28196 142924 28252
rect 142716 28186 142980 28196
rect 142716 26684 142980 26694
rect 142772 26628 142820 26684
rect 142876 26628 142924 26684
rect 142716 26618 142980 26628
rect 142716 25116 142980 25126
rect 142772 25060 142820 25116
rect 142876 25060 142924 25116
rect 142716 25050 142980 25060
rect 142716 23548 142980 23558
rect 142772 23492 142820 23548
rect 142876 23492 142924 23548
rect 142716 23482 142980 23492
rect 142716 21980 142980 21990
rect 142772 21924 142820 21980
rect 142876 21924 142924 21980
rect 142716 21914 142980 21924
rect 142716 20412 142980 20422
rect 142772 20356 142820 20412
rect 142876 20356 142924 20412
rect 142716 20346 142980 20356
rect 142716 18844 142980 18854
rect 142772 18788 142820 18844
rect 142876 18788 142924 18844
rect 142716 18778 142980 18788
rect 145852 17668 145908 17678
rect 142716 17276 142980 17286
rect 142772 17220 142820 17276
rect 142876 17220 142924 17276
rect 142716 17210 142980 17220
rect 142716 15708 142980 15718
rect 142772 15652 142820 15708
rect 142876 15652 142924 15708
rect 142716 15642 142980 15652
rect 142716 14140 142980 14150
rect 142772 14084 142820 14140
rect 142876 14084 142924 14140
rect 142716 14074 142980 14084
rect 143612 12964 143668 12974
rect 142716 12572 142980 12582
rect 142772 12516 142820 12572
rect 142876 12516 142924 12572
rect 142716 12506 142980 12516
rect 142716 11004 142980 11014
rect 142772 10948 142820 11004
rect 142876 10948 142924 11004
rect 142716 10938 142980 10948
rect 142716 9436 142980 9446
rect 142772 9380 142820 9436
rect 142876 9380 142924 9436
rect 142716 9370 142980 9380
rect 141932 9202 141988 9212
rect 142156 8148 142212 8158
rect 142156 8054 142212 8092
rect 143276 8034 143332 8046
rect 143276 7982 143278 8034
rect 143330 7982 143332 8034
rect 142716 7868 142980 7878
rect 142772 7812 142820 7868
rect 142876 7812 142924 7868
rect 142716 7802 142980 7812
rect 142940 7700 142996 7710
rect 142940 7586 142996 7644
rect 143276 7700 143332 7982
rect 143276 7634 143332 7644
rect 142940 7534 142942 7586
rect 142994 7534 142996 7586
rect 141820 7476 141876 7486
rect 141820 7474 141988 7476
rect 141820 7422 141822 7474
rect 141874 7422 141988 7474
rect 141820 7420 141988 7422
rect 141820 7410 141876 7420
rect 141820 6690 141876 6702
rect 141820 6638 141822 6690
rect 141874 6638 141876 6690
rect 141820 6468 141876 6638
rect 141820 6402 141876 6412
rect 141820 5906 141876 5918
rect 141820 5854 141822 5906
rect 141874 5854 141876 5906
rect 141820 5684 141876 5854
rect 141820 5618 141876 5628
rect 141820 5460 141876 5470
rect 141820 5122 141876 5404
rect 141932 5348 141988 7420
rect 142492 6692 142548 6702
rect 142492 6598 142548 6636
rect 142940 6692 142996 7534
rect 142940 6690 143108 6692
rect 142940 6638 142942 6690
rect 142994 6638 143108 6690
rect 142940 6636 143108 6638
rect 142940 6626 142996 6636
rect 142716 6300 142980 6310
rect 142772 6244 142820 6300
rect 142876 6244 142924 6300
rect 142716 6234 142980 6244
rect 141932 5282 141988 5292
rect 142492 5236 142548 5246
rect 141820 5070 141822 5122
rect 141874 5070 141876 5122
rect 141820 5058 141876 5070
rect 142268 5124 142324 5134
rect 141484 4946 141540 4956
rect 141260 4340 141316 4350
rect 141260 3442 141316 4284
rect 142268 4338 142324 5068
rect 142492 5122 142548 5180
rect 142492 5070 142494 5122
rect 142546 5070 142548 5122
rect 142492 5058 142548 5070
rect 143052 5124 143108 6636
rect 143052 5030 143108 5068
rect 142716 4732 142980 4742
rect 142772 4676 142820 4732
rect 142876 4676 142924 4732
rect 142716 4666 142980 4676
rect 142268 4286 142270 4338
rect 142322 4286 142324 4338
rect 142268 4274 142324 4286
rect 143500 4340 143556 4350
rect 143500 4246 143556 4284
rect 143052 4228 143108 4238
rect 143052 4134 143108 4172
rect 142828 3668 142884 3678
rect 142828 3574 142884 3612
rect 143612 3668 143668 12908
rect 144732 8370 144788 8382
rect 144732 8318 144734 8370
rect 144786 8318 144788 8370
rect 144060 8034 144116 8046
rect 144060 7982 144062 8034
rect 144114 7982 144116 8034
rect 144060 7476 144116 7982
rect 144060 7382 144116 7420
rect 144732 6804 144788 8318
rect 145180 8034 145236 8046
rect 145180 7982 145182 8034
rect 145234 7982 145236 8034
rect 145180 7140 145236 7982
rect 145180 7074 145236 7084
rect 145292 8036 145348 8046
rect 145180 6916 145236 6926
rect 145068 6804 145124 6814
rect 144732 6748 145068 6804
rect 144620 6580 144676 6590
rect 144620 6486 144676 6524
rect 144284 6468 144340 6478
rect 144340 6412 144452 6468
rect 144284 6374 144340 6412
rect 143612 3602 143668 3612
rect 143948 5906 144004 5918
rect 143948 5854 143950 5906
rect 144002 5854 144004 5906
rect 141260 3390 141262 3442
rect 141314 3390 141316 3442
rect 141260 3378 141316 3390
rect 143388 3444 143444 3454
rect 143612 3444 143668 3454
rect 143388 3442 143668 3444
rect 143388 3390 143390 3442
rect 143442 3390 143614 3442
rect 143666 3390 143668 3442
rect 143388 3388 143668 3390
rect 142716 3164 142980 3174
rect 142772 3108 142820 3164
rect 142876 3108 142924 3164
rect 142716 3098 142980 3108
rect 141036 2594 141092 2604
rect 143388 800 143444 3388
rect 143612 3378 143668 3388
rect 143948 3442 144004 5854
rect 144284 5684 144340 5694
rect 144284 5122 144340 5628
rect 144284 5070 144286 5122
rect 144338 5070 144340 5122
rect 144284 5058 144340 5070
rect 143948 3390 143950 3442
rect 144002 3390 144004 3442
rect 143948 3378 144004 3390
rect 144396 1652 144452 6412
rect 145068 6018 145124 6748
rect 145068 5966 145070 6018
rect 145122 5966 145124 6018
rect 144956 5124 145012 5134
rect 144956 5030 145012 5068
rect 144956 4452 145012 4462
rect 145068 4452 145124 5966
rect 145180 4562 145236 6860
rect 145292 6130 145348 7980
rect 145740 7700 145796 7710
rect 145740 7474 145796 7644
rect 145740 7422 145742 7474
rect 145794 7422 145796 7474
rect 145404 7140 145460 7150
rect 145404 6690 145460 7084
rect 145404 6638 145406 6690
rect 145458 6638 145460 6690
rect 145404 6626 145460 6638
rect 145292 6078 145294 6130
rect 145346 6078 145348 6130
rect 145292 6066 145348 6078
rect 145740 5572 145796 7422
rect 145852 6692 145908 17612
rect 148204 13524 148260 13534
rect 146412 12852 146468 12862
rect 146300 12796 146412 12852
rect 146188 11170 146244 11182
rect 146188 11118 146190 11170
rect 146242 11118 146244 11170
rect 146188 10500 146244 11118
rect 146188 10434 146244 10444
rect 146076 9492 146132 9502
rect 146076 7474 146132 9436
rect 146076 7422 146078 7474
rect 146130 7422 146132 7474
rect 146076 7410 146132 7422
rect 145852 6598 145908 6636
rect 146300 6468 146356 12796
rect 146412 12786 146468 12796
rect 147756 11732 147812 11742
rect 146860 11508 146916 11518
rect 146860 11414 146916 11452
rect 147308 11508 147364 11518
rect 147308 11414 147364 11452
rect 147532 11394 147588 11406
rect 147532 11342 147534 11394
rect 147586 11342 147588 11394
rect 147532 10500 147588 11342
rect 147532 10406 147588 10444
rect 145740 5506 145796 5516
rect 145852 6412 146356 6468
rect 146412 7474 146468 7486
rect 146412 7422 146414 7474
rect 146466 7422 146468 7474
rect 145404 5460 145460 5470
rect 145404 5236 145460 5404
rect 145180 4510 145182 4562
rect 145234 4510 145236 4562
rect 145180 4498 145236 4510
rect 145292 5234 145460 5236
rect 145292 5182 145406 5234
rect 145458 5182 145460 5234
rect 145292 5180 145460 5182
rect 144956 4450 145124 4452
rect 144956 4398 144958 4450
rect 145010 4398 145124 4450
rect 144956 4396 145124 4398
rect 144956 4386 145012 4396
rect 144508 4228 144564 4238
rect 144508 2212 144564 4172
rect 145292 3388 145348 5180
rect 145404 5170 145460 5180
rect 145852 5236 145908 6412
rect 146076 5906 146132 5918
rect 146076 5854 146078 5906
rect 146130 5854 146132 5906
rect 146076 5796 146132 5854
rect 146412 5908 146468 7422
rect 147644 7474 147700 7486
rect 147644 7422 147646 7474
rect 147698 7422 147700 7474
rect 147644 7028 147700 7422
rect 147644 6962 147700 6972
rect 147644 6692 147700 6702
rect 147756 6692 147812 11676
rect 148204 11394 148260 13468
rect 150332 11732 150388 45948
rect 152124 45332 152180 49200
rect 156156 46004 156212 49200
rect 158076 46284 158340 46294
rect 158132 46228 158180 46284
rect 158236 46228 158284 46284
rect 158076 46218 158340 46228
rect 160188 46004 160244 49200
rect 164220 46004 164276 49200
rect 168252 47012 168308 49200
rect 168252 46956 168756 47012
rect 168700 46450 168756 46956
rect 168700 46398 168702 46450
rect 168754 46398 168756 46450
rect 156156 46002 156436 46004
rect 156156 45950 156158 46002
rect 156210 45950 156436 46002
rect 156156 45948 156436 45950
rect 156156 45938 156212 45948
rect 152796 45890 152852 45902
rect 152796 45838 152798 45890
rect 152850 45838 152852 45890
rect 152796 45668 152852 45838
rect 156380 45890 156436 45948
rect 160188 46002 160692 46004
rect 160188 45950 160190 46002
rect 160242 45950 160692 46002
rect 160188 45948 160692 45950
rect 160188 45938 160244 45948
rect 156380 45838 156382 45890
rect 156434 45838 156436 45890
rect 156380 45826 156436 45838
rect 160636 45890 160692 45948
rect 164220 46002 164724 46004
rect 164220 45950 164222 46002
rect 164274 45950 164724 46002
rect 164220 45948 164724 45950
rect 164220 45938 164276 45948
rect 160636 45838 160638 45890
rect 160690 45838 160692 45890
rect 160636 45826 160692 45838
rect 164668 45890 164724 45948
rect 168700 46002 168756 46398
rect 168700 45950 168702 46002
rect 168754 45950 168756 46002
rect 168700 45938 168756 45950
rect 169484 46450 169540 46462
rect 169484 46398 169486 46450
rect 169538 46398 169540 46450
rect 164668 45838 164670 45890
rect 164722 45838 164724 45890
rect 164668 45826 164724 45838
rect 169484 45890 169540 46398
rect 172284 46004 172340 49200
rect 172508 46004 172564 46014
rect 172284 46002 172564 46004
rect 172284 45950 172510 46002
rect 172562 45950 172564 46002
rect 172284 45948 172564 45950
rect 169484 45838 169486 45890
rect 169538 45838 169540 45890
rect 169484 45826 169540 45838
rect 172508 45892 172564 45948
rect 176316 46002 176372 49200
rect 176316 45950 176318 46002
rect 176370 45950 176372 46002
rect 172508 45826 172564 45836
rect 173292 45892 173348 45902
rect 173292 45798 173348 45836
rect 176316 45892 176372 45950
rect 180236 46004 180292 46014
rect 180348 46004 180404 49200
rect 184380 47012 184436 49200
rect 184044 46956 184436 47012
rect 180236 46002 180964 46004
rect 180236 45950 180238 46002
rect 180290 45950 180964 46002
rect 180236 45948 180964 45950
rect 180236 45938 180292 45948
rect 176316 45826 176372 45836
rect 177100 45892 177156 45902
rect 177100 45798 177156 45836
rect 180908 45890 180964 45948
rect 180908 45838 180910 45890
rect 180962 45838 180964 45890
rect 180908 45826 180964 45838
rect 184044 46002 184100 46956
rect 184044 45950 184046 46002
rect 184098 45950 184100 46002
rect 184044 45892 184100 45950
rect 187852 46004 187908 46014
rect 188412 46004 188468 49200
rect 188796 46284 189060 46294
rect 188852 46228 188900 46284
rect 188956 46228 189004 46284
rect 188796 46218 189060 46228
rect 187852 46002 188468 46004
rect 187852 45950 187854 46002
rect 187906 45950 188468 46002
rect 187852 45948 188468 45950
rect 187852 45938 187908 45948
rect 184044 45826 184100 45836
rect 184828 45892 184884 45902
rect 188412 45892 188468 45948
rect 192444 46004 192500 49200
rect 192444 46002 192724 46004
rect 192444 45950 192446 46002
rect 192498 45950 192724 46002
rect 192444 45948 192724 45950
rect 192444 45938 192500 45948
rect 188636 45892 188692 45902
rect 188412 45890 188692 45892
rect 188412 45838 188638 45890
rect 188690 45838 188692 45890
rect 188412 45836 188692 45838
rect 184828 45798 184884 45836
rect 188636 45826 188692 45836
rect 192668 45890 192724 45948
rect 192668 45838 192670 45890
rect 192722 45838 192724 45890
rect 192668 45826 192724 45838
rect 193116 46002 193172 46014
rect 193116 45950 193118 46002
rect 193170 45950 193172 46002
rect 187292 45780 187348 45790
rect 153244 45668 153300 45678
rect 152796 45666 153300 45668
rect 152796 45614 153246 45666
rect 153298 45614 153300 45666
rect 152796 45612 153300 45614
rect 152124 45266 152180 45276
rect 152348 45106 152404 45118
rect 152348 45054 152350 45106
rect 152402 45054 152404 45106
rect 152124 44996 152180 45006
rect 152348 44996 152404 45054
rect 152180 44940 152404 44996
rect 152124 44902 152180 44940
rect 153244 12740 153300 45612
rect 156716 45666 156772 45678
rect 156716 45614 156718 45666
rect 156770 45614 156772 45666
rect 153356 45332 153412 45342
rect 153356 45238 153412 45276
rect 156716 43708 156772 45614
rect 160412 45666 160468 45678
rect 160412 45614 160414 45666
rect 160466 45614 160468 45666
rect 158076 44716 158340 44726
rect 158132 44660 158180 44716
rect 158236 44660 158284 44716
rect 158076 44650 158340 44660
rect 156716 43652 157556 43708
rect 153244 12674 153300 12684
rect 153692 14308 153748 14318
rect 150332 11666 150388 11676
rect 150780 12628 150836 12638
rect 149212 11508 149268 11518
rect 150444 11508 150500 11518
rect 150668 11508 150724 11518
rect 148204 11342 148206 11394
rect 148258 11342 148260 11394
rect 147868 11170 147924 11182
rect 147868 11118 147870 11170
rect 147922 11118 147924 11170
rect 147868 11060 147924 11118
rect 147868 11004 148148 11060
rect 147868 10836 147924 10874
rect 147868 10770 147924 10780
rect 148092 10612 148148 11004
rect 148204 10836 148260 11342
rect 148764 11396 148820 11406
rect 148764 11394 148932 11396
rect 148764 11342 148766 11394
rect 148818 11342 148932 11394
rect 148764 11340 148932 11342
rect 148764 11330 148820 11340
rect 148260 10780 148372 10836
rect 148204 10770 148260 10780
rect 147868 10556 148148 10612
rect 148204 10610 148260 10622
rect 148204 10558 148206 10610
rect 148258 10558 148260 10610
rect 147868 8372 147924 10556
rect 148204 10500 148260 10558
rect 148204 10434 148260 10444
rect 148204 9940 148260 9950
rect 148316 9940 148372 10780
rect 148764 10498 148820 10510
rect 148764 10446 148766 10498
rect 148818 10446 148820 10498
rect 148204 9938 148596 9940
rect 148204 9886 148206 9938
rect 148258 9886 148596 9938
rect 148204 9884 148596 9886
rect 148204 9874 148260 9884
rect 148540 9826 148596 9884
rect 148540 9774 148542 9826
rect 148594 9774 148596 9826
rect 148540 9762 148596 9774
rect 148764 9828 148820 10446
rect 148764 9762 148820 9772
rect 148876 10276 148932 11340
rect 149212 10610 149268 11452
rect 150220 11506 150668 11508
rect 150220 11454 150446 11506
rect 150498 11454 150668 11506
rect 150220 11452 150668 11454
rect 150108 11282 150164 11294
rect 150108 11230 150110 11282
rect 150162 11230 150164 11282
rect 149660 10612 149716 10622
rect 149212 10558 149214 10610
rect 149266 10558 149268 10610
rect 149212 10546 149268 10558
rect 149548 10556 149660 10612
rect 147868 8278 147924 8316
rect 147980 9604 148036 9614
rect 147868 7700 147924 7710
rect 147868 7606 147924 7644
rect 147196 6690 147812 6692
rect 147196 6638 147646 6690
rect 147698 6638 147812 6690
rect 147196 6636 147812 6638
rect 147980 6690 148036 9548
rect 148652 9604 148708 9614
rect 148652 9510 148708 9548
rect 148428 9268 148484 9278
rect 148428 9174 148484 9212
rect 148540 9156 148596 9166
rect 148540 9062 148596 9100
rect 148540 8372 148596 8382
rect 148540 8278 148596 8316
rect 148764 8372 148820 8382
rect 148876 8372 148932 10220
rect 149548 10052 149604 10556
rect 149660 10518 149716 10556
rect 149324 9996 149604 10052
rect 149324 9156 149380 9996
rect 149324 9044 149380 9100
rect 149548 9828 149604 9838
rect 149324 9042 149492 9044
rect 149324 8990 149326 9042
rect 149378 8990 149492 9042
rect 149324 8988 149492 8990
rect 149324 8978 149380 8988
rect 149436 8708 149492 8988
rect 149548 9042 149604 9772
rect 149772 9826 149828 9838
rect 149772 9774 149774 9826
rect 149826 9774 149828 9826
rect 149772 9268 149828 9774
rect 150108 9828 150164 11230
rect 150108 9762 150164 9772
rect 149772 9202 149828 9212
rect 149996 9602 150052 9614
rect 149996 9550 149998 9602
rect 150050 9550 150052 9602
rect 149548 8990 149550 9042
rect 149602 8990 149604 9042
rect 149548 8978 149604 8990
rect 149660 8932 149716 8942
rect 149660 8838 149716 8876
rect 149436 8652 149940 8708
rect 148764 8370 148932 8372
rect 148764 8318 148766 8370
rect 148818 8318 148932 8370
rect 148764 8316 148932 8318
rect 149884 8370 149940 8652
rect 149884 8318 149886 8370
rect 149938 8318 149940 8370
rect 148764 8306 148820 8316
rect 149884 8306 149940 8318
rect 148204 8034 148260 8046
rect 148204 7982 148206 8034
rect 148258 7982 148260 8034
rect 147980 6638 147982 6690
rect 148034 6638 148036 6690
rect 146748 5908 146804 5918
rect 146412 5906 146804 5908
rect 146412 5854 146750 5906
rect 146802 5854 146804 5906
rect 146412 5852 146804 5854
rect 146076 5730 146132 5740
rect 145852 5142 145908 5180
rect 146636 5124 146692 5852
rect 146748 5842 146804 5852
rect 147196 5906 147252 6636
rect 147644 6626 147700 6636
rect 147980 6626 148036 6638
rect 148092 7586 148148 7598
rect 148092 7534 148094 7586
rect 148146 7534 148148 7586
rect 148092 6804 148148 7534
rect 147196 5854 147198 5906
rect 147250 5854 147252 5906
rect 147196 5842 147252 5854
rect 147308 6466 147364 6478
rect 147308 6414 147310 6466
rect 147362 6414 147364 6466
rect 147308 5908 147364 6414
rect 147308 5236 147364 5852
rect 147196 5180 147364 5236
rect 146076 4338 146132 4350
rect 146076 4286 146078 4338
rect 146130 4286 146132 4338
rect 146076 3668 146132 4286
rect 146636 4338 146692 5068
rect 146636 4286 146638 4338
rect 146690 4286 146692 4338
rect 146636 4274 146692 4286
rect 146748 5122 146804 5134
rect 146748 5070 146750 5122
rect 146802 5070 146804 5122
rect 146076 3602 146132 3612
rect 145964 3444 146020 3454
rect 146412 3444 146468 3454
rect 145964 3442 146468 3444
rect 145964 3390 145966 3442
rect 146018 3390 146414 3442
rect 146466 3390 146468 3442
rect 145964 3388 146468 3390
rect 145292 3332 145460 3388
rect 145964 3378 146020 3388
rect 144508 2146 144564 2156
rect 144396 1586 144452 1596
rect 145404 1428 145460 3332
rect 145404 1362 145460 1372
rect 146076 800 146132 3388
rect 146412 3378 146468 3388
rect 146748 3442 146804 5070
rect 146860 4900 146916 4910
rect 146860 4806 146916 4844
rect 147084 4340 147140 4350
rect 147084 4246 147140 4284
rect 146748 3390 146750 3442
rect 146802 3390 146804 3442
rect 146748 3378 146804 3390
rect 147196 3388 147252 5180
rect 147420 5012 147476 5022
rect 148092 5012 148148 6748
rect 148204 7476 148260 7982
rect 149996 7700 150052 9550
rect 150108 9492 150164 9502
rect 150108 9266 150164 9436
rect 150108 9214 150110 9266
rect 150162 9214 150164 9266
rect 150108 9202 150164 9214
rect 150220 8258 150276 11452
rect 150444 11442 150500 11452
rect 150668 11442 150724 11452
rect 150556 10276 150612 10286
rect 150556 9714 150612 10220
rect 150556 9662 150558 9714
rect 150610 9662 150612 9714
rect 150556 9650 150612 9662
rect 150220 8206 150222 8258
rect 150274 8206 150276 8258
rect 150220 8194 150276 8206
rect 150668 9604 150724 9614
rect 150668 9042 150724 9548
rect 150780 9492 150836 12572
rect 151228 10612 151284 10622
rect 151228 10518 151284 10556
rect 153132 10610 153188 10622
rect 153132 10558 153134 10610
rect 153186 10558 153188 10610
rect 151788 10500 151844 10510
rect 151788 10498 152180 10500
rect 151788 10446 151790 10498
rect 151842 10446 152180 10498
rect 151788 10444 152180 10446
rect 151788 10434 151844 10444
rect 150780 9426 150836 9436
rect 151452 10164 151508 10174
rect 151116 9268 151172 9278
rect 151452 9268 151508 10108
rect 151564 9828 151620 9838
rect 151900 9828 151956 9838
rect 151620 9826 151956 9828
rect 151620 9774 151902 9826
rect 151954 9774 151956 9826
rect 151620 9772 151956 9774
rect 151564 9734 151620 9772
rect 151900 9762 151956 9772
rect 151676 9604 151732 9614
rect 151564 9268 151620 9278
rect 151452 9266 151620 9268
rect 151452 9214 151566 9266
rect 151618 9214 151620 9266
rect 151452 9212 151620 9214
rect 150668 8990 150670 9042
rect 150722 8990 150724 9042
rect 150668 8146 150724 8990
rect 151004 9154 151060 9166
rect 151004 9102 151006 9154
rect 151058 9102 151060 9154
rect 151004 8260 151060 9102
rect 151004 8194 151060 8204
rect 150668 8094 150670 8146
rect 150722 8094 150724 8146
rect 150668 8082 150724 8094
rect 150220 8036 150276 8046
rect 150220 8034 150388 8036
rect 150220 7982 150222 8034
rect 150274 7982 150388 8034
rect 150220 7980 150388 7982
rect 150220 7970 150276 7980
rect 149996 7644 150276 7700
rect 148204 6692 148260 7420
rect 148764 7476 148820 7486
rect 148652 6692 148708 6702
rect 148204 6690 148708 6692
rect 148204 6638 148654 6690
rect 148706 6638 148708 6690
rect 148204 6636 148708 6638
rect 148652 6626 148708 6636
rect 148316 6468 148372 6478
rect 148764 6468 148820 7420
rect 149324 7474 149380 7486
rect 149324 7422 149326 7474
rect 149378 7422 149380 7474
rect 148316 6466 148820 6468
rect 148316 6414 148318 6466
rect 148370 6414 148820 6466
rect 148316 6412 148820 6414
rect 148876 7364 148932 7374
rect 148316 6402 148372 6412
rect 148540 5906 148596 5918
rect 148540 5854 148542 5906
rect 148594 5854 148596 5906
rect 148540 5572 148596 5854
rect 148428 5516 148540 5572
rect 148204 5012 148260 5022
rect 148092 5010 148260 5012
rect 148092 4958 148206 5010
rect 148258 4958 148260 5010
rect 148092 4956 148260 4958
rect 147420 4228 147476 4956
rect 148204 4946 148260 4956
rect 147420 3666 147476 4172
rect 148316 4340 148372 4350
rect 147420 3614 147422 3666
rect 147474 3614 147476 3666
rect 147420 3602 147476 3614
rect 147868 3778 147924 3790
rect 147868 3726 147870 3778
rect 147922 3726 147924 3778
rect 147868 3666 147924 3726
rect 147868 3614 147870 3666
rect 147922 3614 147924 3666
rect 147868 3602 147924 3614
rect 148316 3666 148372 4284
rect 148428 4338 148484 5516
rect 148540 5506 148596 5516
rect 148540 5124 148596 5134
rect 148540 5010 148596 5068
rect 148540 4958 148542 5010
rect 148594 4958 148596 5010
rect 148540 4946 148596 4958
rect 148428 4286 148430 4338
rect 148482 4286 148484 4338
rect 148428 4274 148484 4286
rect 148876 4338 148932 7308
rect 148988 6468 149044 6478
rect 148988 5122 149044 6412
rect 149100 5796 149156 5806
rect 149156 5740 149268 5796
rect 149100 5702 149156 5740
rect 148988 5070 148990 5122
rect 149042 5070 149044 5122
rect 148988 5058 149044 5070
rect 149100 4564 149156 4574
rect 149100 4470 149156 4508
rect 148876 4286 148878 4338
rect 148930 4286 148932 4338
rect 148876 4274 148932 4286
rect 148764 3780 148820 3790
rect 148764 3778 149044 3780
rect 148764 3726 148766 3778
rect 148818 3726 149044 3778
rect 148764 3724 149044 3726
rect 148764 3714 148820 3724
rect 148316 3614 148318 3666
rect 148370 3614 148372 3666
rect 147196 3332 147364 3388
rect 147308 2436 147364 3332
rect 147308 2370 147364 2380
rect 148316 2436 148372 3614
rect 148652 3668 148708 3678
rect 148652 3556 148708 3612
rect 148764 3556 148820 3566
rect 148652 3554 148820 3556
rect 148652 3502 148766 3554
rect 148818 3502 148820 3554
rect 148652 3500 148820 3502
rect 148764 3490 148820 3500
rect 148316 2370 148372 2380
rect 148988 3442 149044 3724
rect 148988 3390 148990 3442
rect 149042 3390 149044 3442
rect 148988 2212 149044 3390
rect 148764 2156 149044 2212
rect 148764 800 148820 2156
rect 149212 1540 149268 5740
rect 149324 3442 149380 7422
rect 150108 7362 150164 7374
rect 150108 7310 150110 7362
rect 150162 7310 150164 7362
rect 149996 7252 150052 7262
rect 149996 6690 150052 7196
rect 150108 7028 150164 7310
rect 150220 7140 150276 7644
rect 150220 7074 150276 7084
rect 150108 6962 150164 6972
rect 149996 6638 149998 6690
rect 150050 6638 150052 6690
rect 149996 6626 150052 6638
rect 150332 6690 150388 7980
rect 151116 7700 151172 9212
rect 151564 9202 151620 9212
rect 151676 8484 151732 9548
rect 152124 9268 152180 10444
rect 152124 9042 152180 9212
rect 152124 8990 152126 9042
rect 152178 8990 152180 9042
rect 152124 8978 152180 8990
rect 152236 10388 152292 10398
rect 151004 7644 151396 7700
rect 150332 6638 150334 6690
rect 150386 6638 150388 6690
rect 149660 6244 149716 6254
rect 149660 6130 149716 6188
rect 149660 6078 149662 6130
rect 149714 6078 149716 6130
rect 149436 5908 149492 5918
rect 149436 5814 149492 5852
rect 149660 4562 149716 6078
rect 149884 6020 149940 6030
rect 149660 4510 149662 4562
rect 149714 4510 149716 4562
rect 149660 4498 149716 4510
rect 149772 5964 149884 6020
rect 149772 4564 149828 5964
rect 149884 5926 149940 5964
rect 150108 5908 150164 5918
rect 149884 4564 149940 4574
rect 149828 4562 149940 4564
rect 149828 4510 149886 4562
rect 149938 4510 149940 4562
rect 149828 4508 149940 4510
rect 149772 4470 149828 4508
rect 149884 4498 149940 4508
rect 150108 4450 150164 5852
rect 150220 5796 150276 5806
rect 150220 5702 150276 5740
rect 150332 5684 150388 6638
rect 150780 7474 150836 7486
rect 150780 7422 150782 7474
rect 150834 7422 150836 7474
rect 150332 5618 150388 5628
rect 150668 5908 150724 5918
rect 150556 5572 150612 5582
rect 150332 5122 150388 5134
rect 150332 5070 150334 5122
rect 150386 5070 150388 5122
rect 150332 4900 150388 5070
rect 150556 5122 150612 5516
rect 150556 5070 150558 5122
rect 150610 5070 150612 5122
rect 150556 5058 150612 5070
rect 150332 4834 150388 4844
rect 150668 4562 150724 5852
rect 150780 5794 150836 7422
rect 150892 7476 150948 7486
rect 150892 7382 150948 7420
rect 150780 5742 150782 5794
rect 150834 5742 150836 5794
rect 150780 4788 150836 5742
rect 150780 4722 150836 4732
rect 151004 4564 151060 7644
rect 151340 7586 151396 7644
rect 151340 7534 151342 7586
rect 151394 7534 151396 7586
rect 151340 7522 151396 7534
rect 151676 7586 151732 8428
rect 152012 8036 152068 8046
rect 151676 7534 151678 7586
rect 151730 7534 151732 7586
rect 151676 7522 151732 7534
rect 151788 8034 152068 8036
rect 151788 7982 152014 8034
rect 152066 7982 152068 8034
rect 151788 7980 152068 7982
rect 151116 7474 151172 7486
rect 151116 7422 151118 7474
rect 151170 7422 151172 7474
rect 151116 7364 151172 7422
rect 151116 7298 151172 7308
rect 151228 7476 151284 7486
rect 151116 6692 151172 6702
rect 151116 6598 151172 6636
rect 151228 5012 151284 7420
rect 151452 7362 151508 7374
rect 151452 7310 151454 7362
rect 151506 7310 151508 7362
rect 151452 6916 151508 7310
rect 151452 6850 151508 6860
rect 151452 6244 151508 6254
rect 151452 6132 151508 6188
rect 151788 6132 151844 7980
rect 152012 7970 152068 7980
rect 151900 7812 151956 7822
rect 152236 7812 152292 10332
rect 153132 10276 153188 10558
rect 153132 10210 153188 10220
rect 153580 10500 153636 10510
rect 153244 9940 153300 9950
rect 152460 9826 152516 9838
rect 152460 9774 152462 9826
rect 152514 9774 152516 9826
rect 152460 9044 152516 9774
rect 152348 8260 152404 8270
rect 152348 8166 152404 8204
rect 152460 7812 152516 8988
rect 152796 8484 152852 8494
rect 152796 8370 152852 8428
rect 152796 8318 152798 8370
rect 152850 8318 152852 8370
rect 152796 8306 152852 8318
rect 153020 8482 153076 8494
rect 153020 8430 153022 8482
rect 153074 8430 153076 8482
rect 151900 7698 151956 7756
rect 151900 7646 151902 7698
rect 151954 7646 151956 7698
rect 151900 7634 151956 7646
rect 152012 7756 152292 7812
rect 152348 7756 152516 7812
rect 151900 6804 151956 6814
rect 152012 6804 152068 7756
rect 152348 7700 152404 7756
rect 152236 7644 152404 7700
rect 152124 7476 152180 7486
rect 152124 7382 152180 7420
rect 152236 7364 152292 7644
rect 152684 7588 152740 7598
rect 152236 7298 152292 7308
rect 152348 7586 152740 7588
rect 152348 7534 152686 7586
rect 152738 7534 152740 7586
rect 152348 7532 152740 7534
rect 152348 7474 152404 7532
rect 152684 7522 152740 7532
rect 152348 7422 152350 7474
rect 152402 7422 152404 7474
rect 151900 6802 152068 6804
rect 151900 6750 151902 6802
rect 151954 6750 152068 6802
rect 151900 6748 152068 6750
rect 152124 7140 152180 7150
rect 151900 6738 151956 6748
rect 152124 6578 152180 7084
rect 152124 6526 152126 6578
rect 152178 6526 152180 6578
rect 152124 6514 152180 6526
rect 151452 6076 151844 6132
rect 151452 6018 151508 6076
rect 151452 5966 151454 6018
rect 151506 5966 151508 6018
rect 151452 5954 151508 5966
rect 151340 5908 151396 5918
rect 151340 5814 151396 5852
rect 151228 4946 151284 4956
rect 151788 4900 151844 6076
rect 152124 6020 152180 6030
rect 151900 5908 151956 5918
rect 151900 5124 151956 5852
rect 152124 5908 152180 5964
rect 152124 5906 152292 5908
rect 152124 5854 152126 5906
rect 152178 5854 152292 5906
rect 152124 5852 152292 5854
rect 152124 5842 152180 5852
rect 152012 5124 152068 5134
rect 151900 5122 152068 5124
rect 151900 5070 152014 5122
rect 152066 5070 152068 5122
rect 151900 5068 152068 5070
rect 152012 5058 152068 5068
rect 152236 5122 152292 5852
rect 152236 5070 152238 5122
rect 152290 5070 152292 5122
rect 152236 5058 152292 5070
rect 151788 4844 152292 4900
rect 150668 4510 150670 4562
rect 150722 4510 150724 4562
rect 150668 4498 150724 4510
rect 150892 4562 151060 4564
rect 150892 4510 151006 4562
rect 151058 4510 151060 4562
rect 150892 4508 151060 4510
rect 150108 4398 150110 4450
rect 150162 4398 150164 4450
rect 150108 4386 150164 4398
rect 150220 4452 150276 4462
rect 150220 4358 150276 4396
rect 149436 4338 149492 4350
rect 149436 4286 149438 4338
rect 149490 4286 149492 4338
rect 149436 4004 149492 4286
rect 149436 3938 149492 3948
rect 150332 4004 150388 4014
rect 150332 3666 150388 3948
rect 150332 3614 150334 3666
rect 150386 3614 150388 3666
rect 150332 3602 150388 3614
rect 150892 3554 150948 4508
rect 151004 4498 151060 4508
rect 151452 4338 151508 4350
rect 151452 4286 151454 4338
rect 151506 4286 151508 4338
rect 150892 3502 150894 3554
rect 150946 3502 150948 3554
rect 150892 3490 150948 3502
rect 151228 4226 151284 4238
rect 151228 4174 151230 4226
rect 151282 4174 151284 4226
rect 149324 3390 149326 3442
rect 149378 3390 149380 3442
rect 149324 3378 149380 3390
rect 151228 2324 151284 4174
rect 151452 3892 151508 4286
rect 151452 3826 151508 3836
rect 152012 3780 152068 3790
rect 151340 3554 151396 3566
rect 151340 3502 151342 3554
rect 151394 3502 151396 3554
rect 151340 3444 151396 3502
rect 151340 3378 151396 3388
rect 151452 3556 151508 3566
rect 151228 2258 151284 2268
rect 149212 1474 149268 1484
rect 151452 800 151508 3500
rect 152012 3554 152068 3724
rect 152012 3502 152014 3554
rect 152066 3502 152068 3554
rect 152012 3490 152068 3502
rect 152236 3554 152292 4844
rect 152348 4452 152404 7422
rect 152908 7476 152964 7486
rect 152908 7382 152964 7420
rect 152460 7364 152516 7374
rect 152460 7270 152516 7308
rect 152796 7250 152852 7262
rect 152796 7198 152798 7250
rect 152850 7198 152852 7250
rect 152684 6356 152740 6366
rect 152572 6244 152628 6254
rect 152460 6132 152516 6142
rect 152460 5906 152516 6076
rect 152460 5854 152462 5906
rect 152514 5854 152516 5906
rect 152460 5842 152516 5854
rect 152572 5346 152628 6188
rect 152684 6018 152740 6300
rect 152684 5966 152686 6018
rect 152738 5966 152740 6018
rect 152684 5954 152740 5966
rect 152572 5294 152574 5346
rect 152626 5294 152628 5346
rect 152572 5282 152628 5294
rect 152796 5236 152852 7198
rect 153020 5908 153076 8430
rect 153244 8484 153300 9884
rect 153356 9156 153412 9166
rect 153580 9156 153636 10444
rect 153356 9154 153636 9156
rect 153356 9102 153358 9154
rect 153410 9102 153636 9154
rect 153356 9100 153636 9102
rect 153356 9090 153412 9100
rect 153132 7812 153188 7822
rect 153132 7698 153188 7756
rect 153132 7646 153134 7698
rect 153186 7646 153188 7698
rect 153132 7634 153188 7646
rect 153244 7474 153300 8428
rect 153468 8820 153524 8830
rect 153244 7422 153246 7474
rect 153298 7422 153300 7474
rect 153244 7410 153300 7422
rect 153356 8034 153412 8046
rect 153356 7982 153358 8034
rect 153410 7982 153412 8034
rect 153356 6916 153412 7982
rect 153244 6860 153412 6916
rect 153244 6468 153300 6860
rect 153244 6402 153300 6412
rect 153356 6690 153412 6702
rect 153356 6638 153358 6690
rect 153410 6638 153412 6690
rect 153020 5852 153300 5908
rect 153132 5684 153188 5694
rect 152796 5170 152852 5180
rect 152908 5682 153188 5684
rect 152908 5630 153134 5682
rect 153186 5630 153188 5682
rect 152908 5628 153188 5630
rect 152572 5122 152628 5134
rect 152572 5070 152574 5122
rect 152626 5070 152628 5122
rect 152460 5012 152516 5022
rect 152460 4918 152516 4956
rect 152572 4676 152628 5070
rect 152572 4610 152628 4620
rect 152796 4452 152852 4462
rect 152348 4450 152852 4452
rect 152348 4398 152798 4450
rect 152850 4398 152852 4450
rect 152348 4396 152852 4398
rect 152236 3502 152238 3554
rect 152290 3502 152292 3554
rect 152236 3490 152292 3502
rect 152460 3892 152516 3902
rect 152460 3554 152516 3836
rect 152460 3502 152462 3554
rect 152514 3502 152516 3554
rect 152460 3490 152516 3502
rect 152684 3554 152740 4396
rect 152796 4386 152852 4396
rect 152796 3668 152852 3678
rect 152796 3574 152852 3612
rect 152684 3502 152686 3554
rect 152738 3502 152740 3554
rect 152572 3444 152628 3454
rect 152684 3444 152740 3502
rect 152628 3388 152740 3444
rect 152572 3378 152628 3388
rect 152908 2548 152964 5628
rect 153132 5618 153188 5628
rect 153020 5348 153076 5358
rect 153020 5254 153076 5292
rect 153244 4900 153300 5852
rect 153244 4834 153300 4844
rect 153356 4676 153412 6638
rect 153468 5122 153524 8764
rect 153580 8372 153636 8382
rect 153692 8372 153748 14252
rect 154588 12740 154644 12750
rect 154028 10724 154084 10734
rect 154028 9602 154084 10668
rect 154588 10498 154644 12684
rect 156492 12178 156548 12190
rect 156492 12126 156494 12178
rect 156546 12126 156548 12178
rect 156044 12066 156100 12078
rect 156044 12014 156046 12066
rect 156098 12014 156100 12066
rect 155260 11564 155764 11620
rect 155260 11506 155316 11564
rect 155260 11454 155262 11506
rect 155314 11454 155316 11506
rect 155260 11442 155316 11454
rect 155596 11394 155652 11406
rect 155596 11342 155598 11394
rect 155650 11342 155652 11394
rect 155148 10948 155204 10958
rect 154924 10724 154980 10734
rect 154924 10630 154980 10668
rect 154588 10446 154590 10498
rect 154642 10446 154644 10498
rect 154588 10434 154644 10446
rect 154812 10276 154868 10286
rect 154812 9826 154868 10220
rect 154812 9774 154814 9826
rect 154866 9774 154868 9826
rect 154812 9762 154868 9774
rect 155148 9714 155204 10892
rect 155596 10500 155652 11342
rect 155596 10434 155652 10444
rect 155708 10610 155764 11564
rect 155708 10558 155710 10610
rect 155762 10558 155764 10610
rect 155596 10052 155652 10062
rect 155596 9826 155652 9996
rect 155596 9774 155598 9826
rect 155650 9774 155652 9826
rect 155596 9762 155652 9774
rect 155148 9662 155150 9714
rect 155202 9662 155204 9714
rect 155148 9650 155204 9662
rect 154028 9550 154030 9602
rect 154082 9550 154084 9602
rect 153916 9044 153972 9054
rect 153580 8370 153748 8372
rect 153580 8318 153582 8370
rect 153634 8318 153694 8370
rect 153746 8318 153748 8370
rect 153580 8316 153748 8318
rect 153580 8306 153636 8316
rect 153692 8306 153748 8316
rect 153804 8484 153860 8494
rect 153804 7698 153860 8428
rect 153804 7646 153806 7698
rect 153858 7646 153860 7698
rect 153804 7634 153860 7646
rect 153468 5070 153470 5122
rect 153522 5070 153524 5122
rect 153468 5058 153524 5070
rect 153580 7476 153636 7486
rect 153020 4620 153412 4676
rect 153020 3442 153076 4620
rect 153580 3892 153636 7420
rect 153916 6804 153972 8988
rect 154028 7364 154084 9550
rect 155708 9604 155764 10558
rect 156044 11396 156100 12014
rect 156492 11508 156548 12126
rect 156492 11442 156548 11452
rect 156604 11618 156660 11630
rect 156604 11566 156606 11618
rect 156658 11566 156660 11618
rect 156044 10610 156100 11340
rect 156492 11284 156548 11294
rect 156268 11282 156548 11284
rect 156268 11230 156494 11282
rect 156546 11230 156548 11282
rect 156268 11228 156548 11230
rect 156156 10724 156212 10734
rect 156268 10724 156324 11228
rect 156492 11218 156548 11228
rect 156156 10722 156324 10724
rect 156156 10670 156158 10722
rect 156210 10670 156324 10722
rect 156156 10668 156324 10670
rect 156156 10658 156212 10668
rect 156044 10558 156046 10610
rect 156098 10558 156100 10610
rect 155932 9828 155988 9838
rect 156044 9828 156100 10558
rect 155932 9826 156044 9828
rect 155932 9774 155934 9826
rect 155986 9774 156044 9826
rect 155932 9772 156044 9774
rect 155932 9762 155988 9772
rect 156044 9734 156100 9772
rect 156156 9828 156212 9838
rect 156268 9828 156324 10668
rect 156156 9826 156268 9828
rect 156156 9774 156158 9826
rect 156210 9774 156268 9826
rect 156156 9772 156268 9774
rect 156324 9772 156548 9828
rect 156156 9762 156212 9772
rect 156268 9762 156324 9772
rect 155372 8484 155428 8494
rect 154700 8036 154756 8046
rect 154588 8034 154756 8036
rect 154588 7982 154702 8034
rect 154754 7982 154756 8034
rect 154588 7980 154756 7982
rect 154252 7364 154308 7374
rect 154588 7364 154644 7980
rect 154700 7970 154756 7980
rect 155148 7700 155204 7710
rect 154812 7364 154868 7374
rect 154028 7362 154644 7364
rect 154028 7310 154254 7362
rect 154306 7310 154644 7362
rect 154028 7308 154644 7310
rect 154700 7362 154868 7364
rect 154700 7310 154814 7362
rect 154866 7310 154868 7362
rect 154700 7308 154868 7310
rect 153804 6748 153972 6804
rect 154252 6916 154308 7308
rect 153692 5908 153748 5918
rect 153692 5122 153748 5852
rect 153692 5070 153694 5122
rect 153746 5070 153748 5122
rect 153692 5058 153748 5070
rect 153692 4450 153748 4462
rect 153692 4398 153694 4450
rect 153746 4398 153748 4450
rect 153692 4228 153748 4398
rect 153692 4162 153748 4172
rect 153580 3826 153636 3836
rect 153356 3556 153412 3566
rect 153804 3556 153860 6748
rect 154028 6466 154084 6478
rect 154028 6414 154030 6466
rect 154082 6414 154084 6466
rect 154028 6132 154084 6414
rect 154028 6066 154084 6076
rect 153916 5906 153972 5918
rect 153916 5854 153918 5906
rect 153970 5854 153972 5906
rect 153916 5460 153972 5854
rect 153916 5394 153972 5404
rect 154140 5908 154196 5918
rect 154252 5908 154308 6860
rect 154700 6692 154756 7308
rect 154812 7298 154868 7308
rect 154924 7364 154980 7374
rect 154980 7308 155092 7364
rect 154924 7298 154980 7308
rect 154700 6356 154756 6636
rect 154700 6300 154868 6356
rect 154140 5906 154308 5908
rect 154140 5854 154142 5906
rect 154194 5854 154308 5906
rect 154140 5852 154308 5854
rect 154700 6018 154756 6030
rect 154700 5966 154702 6018
rect 154754 5966 154756 6018
rect 153916 5236 153972 5246
rect 153972 5180 154084 5236
rect 153916 5170 153972 5180
rect 154028 5122 154084 5180
rect 154028 5070 154030 5122
rect 154082 5070 154084 5122
rect 154028 5058 154084 5070
rect 153916 5010 153972 5022
rect 153916 4958 153918 5010
rect 153970 4958 153972 5010
rect 153916 4564 153972 4958
rect 153916 4498 153972 4508
rect 154140 4228 154196 5852
rect 154588 5124 154644 5134
rect 154700 5124 154756 5966
rect 154812 6020 154868 6300
rect 154812 5954 154868 5964
rect 154588 5122 154700 5124
rect 154588 5070 154590 5122
rect 154642 5070 154700 5122
rect 154588 5068 154700 5070
rect 154588 5058 154644 5068
rect 154700 5030 154756 5068
rect 154924 5460 154980 5470
rect 154812 4900 154868 4910
rect 154812 4806 154868 4844
rect 154924 4900 154980 5404
rect 155036 5124 155092 7308
rect 155148 7362 155204 7644
rect 155148 7310 155150 7362
rect 155202 7310 155204 7362
rect 155148 7252 155204 7310
rect 155148 7186 155204 7196
rect 155372 6802 155428 8428
rect 155372 6750 155374 6802
rect 155426 6750 155428 6802
rect 155372 6738 155428 6750
rect 155596 6692 155652 6702
rect 155708 6692 155764 9548
rect 156268 9602 156324 9614
rect 156268 9550 156270 9602
rect 156322 9550 156324 9602
rect 156268 9492 156324 9550
rect 156156 9436 156324 9492
rect 156044 9268 156100 9278
rect 156044 9174 156100 9212
rect 155596 6690 155764 6692
rect 155596 6638 155598 6690
rect 155650 6638 155764 6690
rect 155596 6636 155764 6638
rect 155820 6916 155876 6926
rect 155820 6690 155876 6860
rect 155820 6638 155822 6690
rect 155874 6638 155876 6690
rect 155596 6626 155652 6636
rect 155820 6626 155876 6638
rect 156044 6468 156100 6478
rect 155932 5794 155988 5806
rect 155932 5742 155934 5794
rect 155986 5742 155988 5794
rect 155932 5460 155988 5742
rect 155932 5394 155988 5404
rect 155148 5348 155204 5358
rect 155820 5348 155876 5358
rect 155148 5346 155652 5348
rect 155148 5294 155150 5346
rect 155202 5294 155652 5346
rect 155148 5292 155652 5294
rect 155148 5282 155204 5292
rect 155372 5124 155428 5134
rect 155036 5122 155428 5124
rect 155036 5070 155374 5122
rect 155426 5070 155428 5122
rect 155036 5068 155428 5070
rect 155372 5058 155428 5068
rect 155596 5122 155652 5292
rect 155596 5070 155598 5122
rect 155650 5070 155652 5122
rect 155596 5058 155652 5070
rect 155708 5292 155820 5348
rect 155708 5122 155764 5292
rect 155820 5282 155876 5292
rect 156044 5236 156100 6412
rect 155932 5180 156100 5236
rect 155708 5070 155710 5122
rect 155762 5070 155764 5122
rect 155708 5058 155764 5070
rect 155820 5124 155876 5134
rect 155036 4900 155092 4910
rect 154924 4898 155428 4900
rect 154924 4846 155038 4898
rect 155090 4846 155428 4898
rect 154924 4844 155428 4846
rect 154924 4676 154980 4844
rect 155036 4834 155092 4844
rect 154588 4620 154980 4676
rect 155036 4676 155092 4686
rect 154588 4338 154644 4620
rect 155036 4562 155092 4620
rect 155036 4510 155038 4562
rect 155090 4510 155092 4562
rect 155036 4498 155092 4510
rect 155260 4564 155316 4574
rect 155260 4470 155316 4508
rect 155372 4562 155428 4844
rect 155372 4510 155374 4562
rect 155426 4510 155428 4562
rect 155372 4498 155428 4510
rect 155820 4450 155876 5068
rect 155820 4398 155822 4450
rect 155874 4398 155876 4450
rect 155820 4386 155876 4398
rect 155596 4340 155652 4350
rect 154588 4286 154590 4338
rect 154642 4286 154644 4338
rect 154588 4274 154644 4286
rect 155484 4338 155652 4340
rect 155484 4286 155598 4338
rect 155650 4286 155652 4338
rect 155484 4284 155652 4286
rect 154140 4162 154196 4172
rect 154476 3892 154532 3902
rect 155484 3892 155540 4284
rect 155596 4274 155652 4284
rect 154476 3666 154532 3836
rect 154476 3614 154478 3666
rect 154530 3614 154532 3666
rect 154476 3602 154532 3614
rect 155260 3836 155540 3892
rect 154028 3556 154084 3566
rect 153804 3554 154084 3556
rect 153804 3502 154030 3554
rect 154082 3502 154084 3554
rect 153804 3500 154084 3502
rect 153356 3462 153412 3500
rect 154028 3490 154084 3500
rect 155036 3554 155092 3566
rect 155036 3502 155038 3554
rect 155090 3502 155092 3554
rect 153020 3390 153022 3442
rect 153074 3390 153076 3442
rect 153020 3378 153076 3390
rect 154140 3444 154196 3454
rect 152908 2482 152964 2492
rect 154140 800 154196 3388
rect 155036 3444 155092 3502
rect 155036 3378 155092 3388
rect 155260 3442 155316 3836
rect 155708 3556 155764 3566
rect 155708 3462 155764 3500
rect 155932 3556 155988 5180
rect 156156 5122 156212 9436
rect 156492 8930 156548 9772
rect 156604 9156 156660 11566
rect 157164 11620 157220 11630
rect 156716 11396 156772 11406
rect 156716 11302 156772 11340
rect 157164 11394 157220 11564
rect 157164 11342 157166 11394
rect 157218 11342 157220 11394
rect 157164 11330 157220 11342
rect 156940 11170 156996 11182
rect 156940 11118 156942 11170
rect 156994 11118 156996 11170
rect 156716 11060 156772 11070
rect 156716 10500 156772 11004
rect 156940 10948 156996 11118
rect 156940 10882 156996 10892
rect 156716 10434 156772 10444
rect 157164 10052 157220 10062
rect 156828 9828 156884 9838
rect 156828 9734 156884 9772
rect 157052 9716 157108 9726
rect 157052 9622 157108 9660
rect 156716 9602 156772 9614
rect 156716 9550 156718 9602
rect 156770 9550 156772 9602
rect 156716 9268 156772 9550
rect 156716 9212 156884 9268
rect 156604 9100 156772 9156
rect 156492 8878 156494 8930
rect 156546 8878 156548 8930
rect 156492 8866 156548 8878
rect 156380 8148 156436 8158
rect 156436 8092 156548 8148
rect 156380 8082 156436 8092
rect 156380 5908 156436 5918
rect 156156 5070 156158 5122
rect 156210 5070 156212 5122
rect 156156 5058 156212 5070
rect 156268 5906 156436 5908
rect 156268 5854 156382 5906
rect 156434 5854 156436 5906
rect 156268 5852 156436 5854
rect 156268 5012 156324 5852
rect 156380 5842 156436 5852
rect 156380 5348 156436 5358
rect 156492 5348 156548 8092
rect 156604 7252 156660 7262
rect 156604 6578 156660 7196
rect 156604 6526 156606 6578
rect 156658 6526 156660 6578
rect 156604 6514 156660 6526
rect 156380 5346 156548 5348
rect 156380 5294 156382 5346
rect 156434 5294 156548 5346
rect 156380 5292 156548 5294
rect 156380 5282 156436 5292
rect 156716 5122 156772 9100
rect 156828 8820 156884 9212
rect 157164 9266 157220 9996
rect 157500 9940 157556 43652
rect 158076 43148 158340 43158
rect 158132 43092 158180 43148
rect 158236 43092 158284 43148
rect 158076 43082 158340 43092
rect 158076 41580 158340 41590
rect 158132 41524 158180 41580
rect 158236 41524 158284 41580
rect 158076 41514 158340 41524
rect 158076 40012 158340 40022
rect 158132 39956 158180 40012
rect 158236 39956 158284 40012
rect 158076 39946 158340 39956
rect 158076 38444 158340 38454
rect 158132 38388 158180 38444
rect 158236 38388 158284 38444
rect 158076 38378 158340 38388
rect 158076 36876 158340 36886
rect 158132 36820 158180 36876
rect 158236 36820 158284 36876
rect 158076 36810 158340 36820
rect 158076 35308 158340 35318
rect 158132 35252 158180 35308
rect 158236 35252 158284 35308
rect 158076 35242 158340 35252
rect 158076 33740 158340 33750
rect 158132 33684 158180 33740
rect 158236 33684 158284 33740
rect 158076 33674 158340 33684
rect 158076 32172 158340 32182
rect 158132 32116 158180 32172
rect 158236 32116 158284 32172
rect 158076 32106 158340 32116
rect 158076 30604 158340 30614
rect 158132 30548 158180 30604
rect 158236 30548 158284 30604
rect 158076 30538 158340 30548
rect 158076 29036 158340 29046
rect 158132 28980 158180 29036
rect 158236 28980 158284 29036
rect 158076 28970 158340 28980
rect 158076 27468 158340 27478
rect 158132 27412 158180 27468
rect 158236 27412 158284 27468
rect 158076 27402 158340 27412
rect 158076 25900 158340 25910
rect 158132 25844 158180 25900
rect 158236 25844 158284 25900
rect 158076 25834 158340 25844
rect 158076 24332 158340 24342
rect 158132 24276 158180 24332
rect 158236 24276 158284 24332
rect 158076 24266 158340 24276
rect 158076 22764 158340 22774
rect 158132 22708 158180 22764
rect 158236 22708 158284 22764
rect 158076 22698 158340 22708
rect 158076 21196 158340 21206
rect 158132 21140 158180 21196
rect 158236 21140 158284 21196
rect 158076 21130 158340 21140
rect 158076 19628 158340 19638
rect 158132 19572 158180 19628
rect 158236 19572 158284 19628
rect 158076 19562 158340 19572
rect 158076 18060 158340 18070
rect 158132 18004 158180 18060
rect 158236 18004 158284 18060
rect 158076 17994 158340 18004
rect 158076 16492 158340 16502
rect 158132 16436 158180 16492
rect 158236 16436 158284 16492
rect 158076 16426 158340 16436
rect 158076 14924 158340 14934
rect 158132 14868 158180 14924
rect 158236 14868 158284 14924
rect 158076 14858 158340 14868
rect 158076 13356 158340 13366
rect 158132 13300 158180 13356
rect 158236 13300 158284 13356
rect 158076 13290 158340 13300
rect 158076 11788 158340 11798
rect 158132 11732 158180 11788
rect 158236 11732 158284 11788
rect 158076 11722 158340 11732
rect 157724 11620 157780 11630
rect 157724 11506 157780 11564
rect 157724 11454 157726 11506
rect 157778 11454 157780 11506
rect 157724 11442 157780 11454
rect 160300 11508 160356 11518
rect 159852 11172 159908 11182
rect 158076 10220 158340 10230
rect 158132 10164 158180 10220
rect 158236 10164 158284 10220
rect 158076 10154 158340 10164
rect 157948 9940 158004 9950
rect 157500 9938 158004 9940
rect 157500 9886 157950 9938
rect 158002 9886 158004 9938
rect 157500 9884 158004 9886
rect 157500 9826 157556 9884
rect 157948 9874 158004 9884
rect 157500 9774 157502 9826
rect 157554 9774 157556 9826
rect 157500 9762 157556 9774
rect 157276 9604 157332 9614
rect 157276 9510 157332 9548
rect 157164 9214 157166 9266
rect 157218 9214 157220 9266
rect 157164 9202 157220 9214
rect 156828 8754 156884 8764
rect 158076 8652 158340 8662
rect 158132 8596 158180 8652
rect 158236 8596 158284 8652
rect 158076 8586 158340 8596
rect 156828 8372 156884 8382
rect 156828 6132 156884 8316
rect 159292 8260 159348 8270
rect 158076 7084 158340 7094
rect 158132 7028 158180 7084
rect 158236 7028 158284 7084
rect 158076 7018 158340 7028
rect 156828 6038 156884 6076
rect 157948 6132 158004 6142
rect 157948 6038 158004 6076
rect 159292 6130 159348 8204
rect 159628 6692 159684 6702
rect 159684 6636 159796 6692
rect 159628 6626 159684 6636
rect 159292 6078 159294 6130
rect 159346 6078 159348 6130
rect 157724 6020 157780 6030
rect 157388 5794 157444 5806
rect 157388 5742 157390 5794
rect 157442 5742 157444 5794
rect 157164 5684 157220 5694
rect 156716 5070 156718 5122
rect 156770 5070 156772 5122
rect 156716 5058 156772 5070
rect 156828 5348 156884 5358
rect 156828 5124 156884 5292
rect 156828 5058 156884 5068
rect 157164 5122 157220 5628
rect 157388 5348 157444 5742
rect 157388 5282 157444 5292
rect 157164 5070 157166 5122
rect 157218 5070 157220 5122
rect 157164 5058 157220 5070
rect 157276 5236 157332 5246
rect 157276 5122 157332 5180
rect 157276 5070 157278 5122
rect 157330 5070 157332 5122
rect 157276 5058 157332 5070
rect 157388 5122 157444 5134
rect 157388 5070 157390 5122
rect 157442 5070 157444 5122
rect 156268 4338 156324 4956
rect 156604 5012 156660 5022
rect 156492 4898 156548 4910
rect 156492 4846 156494 4898
rect 156546 4846 156548 4898
rect 156492 4676 156548 4846
rect 156268 4286 156270 4338
rect 156322 4286 156324 4338
rect 156268 4274 156324 4286
rect 156380 4620 156548 4676
rect 156044 3780 156100 3790
rect 156100 3724 156212 3780
rect 156044 3714 156100 3724
rect 156156 3666 156212 3724
rect 156156 3614 156158 3666
rect 156210 3614 156212 3666
rect 156156 3602 156212 3614
rect 155932 3490 155988 3500
rect 155260 3390 155262 3442
rect 155314 3390 155316 3442
rect 155260 3378 155316 3390
rect 156380 2660 156436 4620
rect 156492 4452 156548 4462
rect 156604 4452 156660 4956
rect 156492 4450 156660 4452
rect 156492 4398 156494 4450
rect 156546 4398 156660 4450
rect 156492 4396 156660 4398
rect 156492 4386 156548 4396
rect 157388 3780 157444 5070
rect 157724 4788 157780 5964
rect 158076 5516 158340 5526
rect 158132 5460 158180 5516
rect 158236 5460 158284 5516
rect 158076 5450 158340 5460
rect 157836 5348 157892 5358
rect 157836 5122 157892 5292
rect 157948 5236 158004 5246
rect 157948 5142 158004 5180
rect 157836 5070 157838 5122
rect 157890 5070 157892 5122
rect 157836 5058 157892 5070
rect 159292 5124 159348 6078
rect 159628 6468 159684 6478
rect 159628 6130 159684 6412
rect 159628 6078 159630 6130
rect 159682 6078 159684 6130
rect 159628 6066 159684 6078
rect 159740 5572 159796 6636
rect 159852 6130 159908 11116
rect 160076 10610 160132 10622
rect 160076 10558 160078 10610
rect 160130 10558 160132 10610
rect 160076 9492 160132 10558
rect 160300 10612 160356 11452
rect 160300 10518 160356 10556
rect 160076 9426 160132 9436
rect 160188 10386 160244 10398
rect 160188 10334 160190 10386
rect 160242 10334 160244 10386
rect 160076 7812 160132 7822
rect 160076 6580 160132 7756
rect 159852 6078 159854 6130
rect 159906 6078 159908 6130
rect 159852 6066 159908 6078
rect 159964 6466 160020 6478
rect 159964 6414 159966 6466
rect 160018 6414 160020 6466
rect 159964 6132 160020 6414
rect 159964 6066 160020 6076
rect 160076 5684 160132 6524
rect 160188 5906 160244 10334
rect 160412 10164 160468 45614
rect 164444 45666 164500 45678
rect 164444 45614 164446 45666
rect 164498 45614 164500 45666
rect 162876 15988 162932 15998
rect 160748 11732 160804 11742
rect 160524 10724 160580 10734
rect 160524 10630 160580 10668
rect 160748 10724 160804 11676
rect 162876 11732 162932 15932
rect 163324 12068 163380 12078
rect 162876 11666 162932 11676
rect 163100 12012 163324 12068
rect 162540 11620 162596 11630
rect 162988 11620 163044 11630
rect 162540 11618 162820 11620
rect 162540 11566 162542 11618
rect 162594 11566 162820 11618
rect 162540 11564 162820 11566
rect 162540 11554 162596 11564
rect 162428 11396 162484 11406
rect 162204 11394 162484 11396
rect 162204 11342 162430 11394
rect 162482 11342 162484 11394
rect 162204 11340 162484 11342
rect 161980 10948 162036 10958
rect 161532 10836 161588 10846
rect 161532 10742 161588 10780
rect 160748 10722 161140 10724
rect 160748 10670 160750 10722
rect 160802 10670 161140 10722
rect 160748 10668 161140 10670
rect 160748 10658 160804 10668
rect 160412 10098 160468 10108
rect 161084 9938 161140 10668
rect 161196 10612 161252 10622
rect 161196 10518 161252 10556
rect 161980 10610 162036 10892
rect 162092 10724 162148 10734
rect 162092 10630 162148 10668
rect 161980 10558 161982 10610
rect 162034 10558 162036 10610
rect 161980 10546 162036 10558
rect 161644 10500 161700 10510
rect 161700 10444 161812 10500
rect 161644 10434 161700 10444
rect 161084 9886 161086 9938
rect 161138 9886 161140 9938
rect 161084 9874 161140 9886
rect 161532 9714 161588 9726
rect 161532 9662 161534 9714
rect 161586 9662 161588 9714
rect 161532 9492 161588 9662
rect 161532 9426 161588 9436
rect 160636 8932 160692 8942
rect 160636 7700 160692 8876
rect 161196 8484 161252 8494
rect 160636 7698 160916 7700
rect 160636 7646 160638 7698
rect 160690 7646 160916 7698
rect 160636 7644 160916 7646
rect 160636 7634 160692 7644
rect 160300 7364 160356 7374
rect 160300 6578 160356 7308
rect 160524 6804 160580 6814
rect 160300 6526 160302 6578
rect 160354 6526 160356 6578
rect 160300 6132 160356 6526
rect 160300 6066 160356 6076
rect 160412 6748 160524 6804
rect 160412 6018 160468 6748
rect 160524 6738 160580 6748
rect 160636 6802 160692 6814
rect 160636 6750 160638 6802
rect 160690 6750 160692 6802
rect 160412 5966 160414 6018
rect 160466 5966 160468 6018
rect 160412 5954 160468 5966
rect 160524 6466 160580 6478
rect 160524 6414 160526 6466
rect 160578 6414 160580 6466
rect 160188 5854 160190 5906
rect 160242 5854 160244 5906
rect 160188 5842 160244 5854
rect 160076 5628 160356 5684
rect 159740 5506 159796 5516
rect 159292 5058 159348 5068
rect 158284 5012 158340 5022
rect 158284 4918 158340 4956
rect 160300 5010 160356 5628
rect 160524 5348 160580 6414
rect 160636 6018 160692 6750
rect 160860 6804 160916 7644
rect 161084 7364 161140 7374
rect 161084 7270 161140 7308
rect 161196 7028 161252 8428
rect 161756 8372 161812 10444
rect 161868 9716 161924 9726
rect 162204 9716 162260 11340
rect 162428 11330 162484 11340
rect 162652 11172 162708 11182
rect 162540 11116 162652 11172
rect 162316 10836 162372 10846
rect 162540 10836 162596 11116
rect 162652 11078 162708 11116
rect 162372 10780 162596 10836
rect 162316 10742 162372 10780
rect 162540 10612 162596 10622
rect 162540 9716 162596 10556
rect 161868 9714 162596 9716
rect 161868 9662 161870 9714
rect 161922 9662 162596 9714
rect 161868 9660 162596 9662
rect 162652 10498 162708 10510
rect 162652 10446 162654 10498
rect 162706 10446 162708 10498
rect 161868 9650 161924 9660
rect 161756 8316 162372 8372
rect 161756 7588 161812 7598
rect 161756 7494 161812 7532
rect 162204 7588 162260 7598
rect 161420 7474 161476 7486
rect 161420 7422 161422 7474
rect 161474 7422 161476 7474
rect 161420 7364 161476 7422
rect 161420 7298 161476 7308
rect 162204 7474 162260 7532
rect 162204 7422 162206 7474
rect 162258 7422 162260 7474
rect 161644 7252 161700 7262
rect 161700 7196 161812 7252
rect 161644 7186 161700 7196
rect 161084 6972 161252 7028
rect 160860 6748 161028 6804
rect 160972 6692 161028 6748
rect 160972 6598 161028 6636
rect 160748 6468 160804 6478
rect 160748 6132 160804 6412
rect 160748 6066 160804 6076
rect 160636 5966 160638 6018
rect 160690 5966 160692 6018
rect 160636 5954 160692 5966
rect 160748 5906 160804 5918
rect 160748 5854 160750 5906
rect 160802 5854 160804 5906
rect 160748 5572 160804 5854
rect 160748 5506 160804 5516
rect 160524 5292 160692 5348
rect 160524 5124 160580 5134
rect 160524 5030 160580 5068
rect 160300 4958 160302 5010
rect 160354 4958 160356 5010
rect 160300 4946 160356 4958
rect 157724 4722 157780 4732
rect 157836 4900 157892 4910
rect 157388 3714 157444 3724
rect 156604 3444 156660 3482
rect 156604 3378 156660 3388
rect 157388 3444 157444 3482
rect 156380 2594 156436 2604
rect 157388 2212 157444 3388
rect 157836 3442 157892 4844
rect 158060 4900 158116 4910
rect 158060 4806 158116 4844
rect 159740 4900 159796 4910
rect 158076 3948 158340 3958
rect 158132 3892 158180 3948
rect 158236 3892 158284 3948
rect 158076 3882 158340 3892
rect 157836 3390 157838 3442
rect 157890 3390 157892 3442
rect 157836 3378 157892 3390
rect 158172 3444 158228 3482
rect 158172 3378 158228 3388
rect 159516 3444 159572 3482
rect 156828 2156 157444 2212
rect 156828 800 156884 2156
rect 159516 800 159572 3388
rect 159740 3330 159796 4844
rect 160636 3780 160692 5292
rect 161084 5122 161140 6972
rect 161532 6804 161588 6814
rect 161532 6710 161588 6748
rect 161084 5070 161086 5122
rect 161138 5070 161140 5122
rect 161084 5058 161140 5070
rect 161196 6692 161252 6702
rect 161196 6130 161252 6636
rect 161420 6580 161476 6590
rect 161420 6486 161476 6524
rect 161644 6468 161700 6478
rect 161644 6374 161700 6412
rect 161196 6078 161198 6130
rect 161250 6078 161252 6130
rect 160860 4900 160916 4910
rect 160636 3714 160692 3724
rect 160748 4898 160916 4900
rect 160748 4846 160862 4898
rect 160914 4846 160916 4898
rect 160748 4844 160916 4846
rect 160076 3444 160132 3482
rect 160076 3378 160132 3388
rect 159740 3278 159742 3330
rect 159794 3278 159796 3330
rect 159740 3266 159796 3278
rect 160748 2772 160804 4844
rect 160860 4834 160916 4844
rect 161196 4788 161252 6078
rect 161756 5906 161812 7196
rect 161756 5854 161758 5906
rect 161810 5854 161812 5906
rect 161756 5460 161812 5854
rect 161980 6356 162036 6366
rect 161756 5394 161812 5404
rect 161868 5796 161924 5806
rect 161868 5234 161924 5740
rect 161868 5182 161870 5234
rect 161922 5182 161924 5234
rect 161868 5170 161924 5182
rect 161980 5236 162036 6300
rect 161980 5170 162036 5180
rect 161532 5124 161588 5134
rect 161532 5030 161588 5068
rect 161756 5010 161812 5022
rect 161756 4958 161758 5010
rect 161810 4958 161812 5010
rect 161420 4900 161476 4910
rect 160972 4732 161364 4788
rect 160860 4564 160916 4574
rect 160972 4564 161028 4732
rect 160860 4562 161028 4564
rect 160860 4510 160862 4562
rect 160914 4510 161028 4562
rect 160860 4508 161028 4510
rect 160860 4498 160916 4508
rect 161308 3780 161364 4732
rect 161420 4562 161476 4844
rect 161420 4510 161422 4562
rect 161474 4510 161476 4562
rect 161420 4498 161476 4510
rect 161756 4564 161812 4958
rect 161756 4498 161812 4508
rect 161980 4676 162036 4686
rect 162204 4676 162260 7422
rect 162316 6130 162372 8316
rect 162428 8260 162484 8270
rect 162428 8166 162484 8204
rect 162540 7476 162596 7486
rect 162540 7382 162596 7420
rect 162652 7140 162708 10446
rect 162764 8596 162820 11564
rect 162876 11170 162932 11182
rect 162876 11118 162878 11170
rect 162930 11118 162932 11170
rect 162876 11060 162932 11118
rect 162876 10994 162932 11004
rect 162988 10948 163044 11564
rect 163100 11394 163156 12012
rect 163324 11974 163380 12012
rect 164444 11844 164500 45614
rect 169260 45666 169316 45678
rect 169260 45614 169262 45666
rect 169314 45614 169316 45666
rect 167132 43764 167188 43774
rect 164444 11778 164500 11788
rect 164668 14196 164724 14206
rect 164668 11506 164724 14140
rect 164668 11454 164670 11506
rect 164722 11454 164724 11506
rect 163100 11342 163102 11394
rect 163154 11342 163156 11394
rect 163100 11330 163156 11342
rect 163996 11396 164052 11406
rect 163996 11302 164052 11340
rect 164668 11396 164724 11454
rect 164668 11330 164724 11340
rect 163436 11282 163492 11294
rect 163436 11230 163438 11282
rect 163490 11230 163492 11282
rect 163324 11172 163380 11182
rect 162988 10834 163044 10892
rect 162988 10782 162990 10834
rect 163042 10782 163044 10834
rect 162988 10770 163044 10782
rect 163212 11170 163380 11172
rect 163212 11118 163326 11170
rect 163378 11118 163380 11170
rect 163212 11116 163380 11118
rect 162764 8530 162820 8540
rect 162764 8036 162820 8046
rect 162764 7942 162820 7980
rect 163212 7700 163268 11116
rect 163324 11106 163380 11116
rect 163324 10612 163380 10622
rect 163436 10612 163492 11230
rect 163548 11172 163604 11182
rect 163660 11172 163716 11182
rect 163884 11172 163940 11182
rect 163604 11170 163716 11172
rect 163604 11118 163662 11170
rect 163714 11118 163716 11170
rect 163604 11116 163716 11118
rect 163548 10834 163604 11116
rect 163660 11106 163716 11116
rect 163772 11170 163940 11172
rect 163772 11118 163886 11170
rect 163938 11118 163940 11170
rect 163772 11116 163940 11118
rect 163548 10782 163550 10834
rect 163602 10782 163604 10834
rect 163548 10770 163604 10782
rect 163772 11060 163828 11116
rect 163884 11106 163940 11116
rect 163772 10834 163828 11004
rect 163772 10782 163774 10834
rect 163826 10782 163828 10834
rect 163772 10770 163828 10782
rect 163996 10836 164052 10846
rect 163996 10722 164052 10780
rect 164444 10836 164500 10846
rect 164444 10742 164500 10780
rect 167132 10836 167188 43708
rect 168028 14420 168084 14430
rect 168028 11732 168084 14364
rect 169260 14196 169316 45614
rect 173068 45666 173124 45678
rect 173068 45614 173070 45666
rect 173122 45614 173124 45666
rect 173068 43764 173124 45614
rect 176876 45666 176932 45678
rect 176876 45614 176878 45666
rect 176930 45614 176932 45666
rect 173436 45500 173700 45510
rect 173492 45444 173540 45500
rect 173596 45444 173644 45500
rect 173436 45434 173700 45444
rect 173436 43932 173700 43942
rect 173492 43876 173540 43932
rect 173596 43876 173644 43932
rect 173436 43866 173700 43876
rect 173068 43698 173124 43708
rect 173436 42364 173700 42374
rect 173492 42308 173540 42364
rect 173596 42308 173644 42364
rect 173436 42298 173700 42308
rect 173436 40796 173700 40806
rect 173492 40740 173540 40796
rect 173596 40740 173644 40796
rect 173436 40730 173700 40740
rect 173436 39228 173700 39238
rect 173492 39172 173540 39228
rect 173596 39172 173644 39228
rect 173436 39162 173700 39172
rect 173436 37660 173700 37670
rect 173492 37604 173540 37660
rect 173596 37604 173644 37660
rect 173436 37594 173700 37604
rect 173436 36092 173700 36102
rect 173492 36036 173540 36092
rect 173596 36036 173644 36092
rect 173436 36026 173700 36036
rect 173436 34524 173700 34534
rect 173492 34468 173540 34524
rect 173596 34468 173644 34524
rect 173436 34458 173700 34468
rect 173436 32956 173700 32966
rect 173492 32900 173540 32956
rect 173596 32900 173644 32956
rect 173436 32890 173700 32900
rect 173436 31388 173700 31398
rect 173492 31332 173540 31388
rect 173596 31332 173644 31388
rect 173436 31322 173700 31332
rect 173436 29820 173700 29830
rect 173492 29764 173540 29820
rect 173596 29764 173644 29820
rect 173436 29754 173700 29764
rect 173436 28252 173700 28262
rect 173492 28196 173540 28252
rect 173596 28196 173644 28252
rect 173436 28186 173700 28196
rect 173436 26684 173700 26694
rect 173492 26628 173540 26684
rect 173596 26628 173644 26684
rect 173436 26618 173700 26628
rect 173436 25116 173700 25126
rect 173492 25060 173540 25116
rect 173596 25060 173644 25116
rect 173436 25050 173700 25060
rect 173436 23548 173700 23558
rect 173492 23492 173540 23548
rect 173596 23492 173644 23548
rect 173436 23482 173700 23492
rect 173436 21980 173700 21990
rect 173492 21924 173540 21980
rect 173596 21924 173644 21980
rect 173436 21914 173700 21924
rect 173436 20412 173700 20422
rect 173492 20356 173540 20412
rect 173596 20356 173644 20412
rect 173436 20346 173700 20356
rect 173436 18844 173700 18854
rect 173492 18788 173540 18844
rect 173596 18788 173644 18844
rect 173436 18778 173700 18788
rect 173436 17276 173700 17286
rect 173492 17220 173540 17276
rect 173596 17220 173644 17276
rect 173436 17210 173700 17220
rect 173436 15708 173700 15718
rect 173492 15652 173540 15708
rect 173596 15652 173644 15708
rect 173436 15642 173700 15652
rect 169260 14130 169316 14140
rect 173436 14140 173700 14150
rect 173492 14084 173540 14140
rect 173596 14084 173644 14140
rect 173436 14074 173700 14084
rect 173436 12572 173700 12582
rect 173492 12516 173540 12572
rect 173596 12516 173644 12572
rect 173436 12506 173700 12516
rect 176876 12068 176932 45614
rect 180684 45666 180740 45678
rect 180684 45614 180686 45666
rect 180738 45614 180740 45666
rect 180684 14420 180740 45614
rect 184604 45666 184660 45678
rect 184604 45614 184606 45666
rect 184658 45614 184660 45666
rect 180684 14354 180740 14364
rect 182252 45556 182308 45566
rect 176876 12002 176932 12012
rect 168028 11666 168084 11676
rect 173436 11004 173700 11014
rect 173492 10948 173540 11004
rect 173596 10948 173644 11004
rect 173436 10938 173700 10948
rect 167132 10770 167188 10780
rect 163996 10670 163998 10722
rect 164050 10670 164052 10722
rect 163996 10658 164052 10670
rect 163380 10556 163492 10612
rect 163324 10518 163380 10556
rect 163436 10386 163492 10398
rect 163436 10334 163438 10386
rect 163490 10334 163492 10386
rect 163436 8484 163492 10334
rect 173436 9436 173700 9446
rect 173492 9380 173540 9436
rect 173596 9380 173644 9436
rect 173436 9370 173700 9380
rect 163436 8418 163492 8428
rect 163996 8596 164052 8606
rect 163212 7644 163492 7700
rect 162652 7074 162708 7084
rect 162764 7586 162820 7598
rect 162764 7534 162766 7586
rect 162818 7534 162820 7586
rect 162316 6078 162318 6130
rect 162370 6078 162372 6130
rect 162316 6066 162372 6078
rect 162428 7028 162484 7038
rect 162428 5908 162484 6972
rect 162764 7028 162820 7534
rect 162988 7588 163044 7598
rect 162988 7474 163044 7532
rect 162988 7422 162990 7474
rect 163042 7422 163044 7474
rect 162988 7410 163044 7422
rect 163324 7474 163380 7486
rect 163324 7422 163326 7474
rect 163378 7422 163380 7474
rect 162876 7252 162932 7262
rect 162876 7250 163268 7252
rect 162876 7198 162878 7250
rect 162930 7198 163268 7250
rect 162876 7196 163268 7198
rect 162876 7186 162932 7196
rect 162764 6962 162820 6972
rect 162764 6804 162820 6814
rect 162764 6802 163044 6804
rect 162764 6750 162766 6802
rect 162818 6750 163044 6802
rect 162764 6748 163044 6750
rect 162764 6738 162820 6748
rect 162652 6692 162708 6730
rect 162652 6626 162708 6636
rect 162876 6580 162932 6590
rect 162876 6486 162932 6524
rect 162764 6132 162820 6142
rect 162540 5908 162596 5918
rect 162428 5906 162596 5908
rect 162428 5854 162542 5906
rect 162594 5854 162596 5906
rect 162428 5852 162596 5854
rect 162540 5842 162596 5852
rect 162316 5460 162372 5470
rect 162316 5122 162372 5404
rect 162316 5070 162318 5122
rect 162370 5070 162372 5122
rect 162316 5058 162372 5070
rect 162764 5122 162820 6076
rect 162988 6018 163044 6748
rect 162988 5966 162990 6018
rect 163042 5966 163044 6018
rect 162988 5954 163044 5966
rect 163100 6580 163156 6590
rect 163100 6466 163156 6524
rect 163100 6414 163102 6466
rect 163154 6414 163156 6466
rect 162876 5348 162932 5358
rect 162876 5234 162932 5292
rect 162876 5182 162878 5234
rect 162930 5182 162932 5234
rect 162876 5170 162932 5182
rect 163100 5348 163156 6414
rect 163212 6018 163268 7196
rect 163324 6804 163380 7422
rect 163324 6738 163380 6748
rect 163212 5966 163214 6018
rect 163266 5966 163268 6018
rect 163212 5954 163268 5966
rect 163324 6244 163380 6254
rect 163324 5906 163380 6188
rect 163324 5854 163326 5906
rect 163378 5854 163380 5906
rect 163324 5842 163380 5854
rect 162764 5070 162766 5122
rect 162818 5070 162820 5122
rect 162764 5058 162820 5070
rect 162988 5012 163044 5022
rect 162988 4918 163044 4956
rect 163100 4676 163156 5292
rect 163324 5236 163380 5246
rect 163324 5122 163380 5180
rect 163324 5070 163326 5122
rect 163378 5070 163380 5122
rect 163324 5058 163380 5070
rect 162036 4620 162260 4676
rect 162988 4620 163156 4676
rect 161644 4338 161700 4350
rect 161644 4286 161646 4338
rect 161698 4286 161700 4338
rect 161644 3892 161700 4286
rect 161980 4338 162036 4620
rect 162988 4564 163044 4620
rect 162876 4508 163044 4564
rect 161980 4286 161982 4338
rect 162034 4286 162036 4338
rect 161980 4274 162036 4286
rect 162204 4452 162260 4462
rect 162204 4338 162260 4396
rect 162764 4452 162820 4462
rect 162764 4358 162820 4396
rect 162204 4286 162206 4338
rect 162258 4286 162260 4338
rect 162204 4274 162260 4286
rect 162428 4338 162484 4350
rect 162428 4286 162430 4338
rect 162482 4286 162484 4338
rect 161756 4116 161812 4126
rect 162428 4116 162484 4286
rect 161756 4114 162484 4116
rect 161756 4062 161758 4114
rect 161810 4062 162484 4114
rect 161756 4060 162484 4062
rect 162876 4116 162932 4508
rect 162988 4340 163044 4350
rect 163436 4340 163492 7644
rect 163548 7586 163604 7598
rect 163548 7534 163550 7586
rect 163602 7534 163604 7586
rect 163548 6132 163604 7534
rect 163548 6066 163604 6076
rect 163660 7250 163716 7262
rect 163660 7198 163662 7250
rect 163714 7198 163716 7250
rect 163548 5906 163604 5918
rect 163548 5854 163550 5906
rect 163602 5854 163604 5906
rect 163548 5460 163604 5854
rect 163548 5394 163604 5404
rect 163660 5122 163716 7198
rect 163884 6690 163940 6702
rect 163884 6638 163886 6690
rect 163938 6638 163940 6690
rect 163884 6580 163940 6638
rect 163884 6514 163940 6524
rect 163772 6468 163828 6478
rect 163772 5796 163828 6412
rect 163996 6468 164052 8540
rect 164332 8036 164388 8046
rect 164108 7364 164164 7374
rect 164108 7362 164276 7364
rect 164108 7310 164110 7362
rect 164162 7310 164276 7362
rect 164108 7308 164276 7310
rect 164108 7298 164164 7308
rect 163996 6402 164052 6412
rect 164220 6692 164276 7308
rect 164220 6132 164276 6636
rect 164332 6692 164388 7980
rect 173436 7868 173700 7878
rect 173492 7812 173540 7868
rect 173596 7812 173644 7868
rect 173436 7802 173700 7812
rect 170492 7364 170548 7374
rect 167804 6804 167860 6814
rect 164332 6690 164948 6692
rect 164332 6638 164334 6690
rect 164386 6638 164948 6690
rect 164332 6636 164948 6638
rect 164332 6626 164388 6636
rect 164444 6466 164500 6478
rect 164444 6414 164446 6466
rect 164498 6414 164500 6466
rect 164444 6244 164500 6414
rect 164556 6468 164612 6478
rect 164556 6374 164612 6412
rect 164444 6188 164612 6244
rect 164220 6066 164276 6076
rect 163996 6020 164052 6030
rect 163996 5926 164052 5964
rect 164108 5908 164164 5918
rect 164108 5814 164164 5852
rect 164220 5908 164276 5918
rect 164220 5906 164388 5908
rect 164220 5854 164222 5906
rect 164274 5854 164388 5906
rect 164220 5852 164388 5854
rect 164220 5842 164276 5852
rect 163772 5730 163828 5740
rect 163660 5070 163662 5122
rect 163714 5070 163716 5122
rect 163660 5058 163716 5070
rect 163772 5572 163828 5582
rect 163772 5122 163828 5516
rect 163772 5070 163774 5122
rect 163826 5070 163828 5122
rect 163772 5058 163828 5070
rect 163996 5236 164052 5246
rect 163996 5122 164052 5180
rect 163996 5070 163998 5122
rect 164050 5070 164052 5122
rect 163996 5058 164052 5070
rect 163772 4900 163828 4910
rect 163660 4564 163716 4574
rect 163660 4470 163716 4508
rect 163772 4562 163828 4844
rect 163772 4510 163774 4562
rect 163826 4510 163828 4562
rect 163772 4498 163828 4510
rect 164220 4676 164276 4686
rect 164220 4450 164276 4620
rect 164220 4398 164222 4450
rect 164274 4398 164276 4450
rect 164220 4386 164276 4398
rect 162988 4338 163492 4340
rect 162988 4286 162990 4338
rect 163042 4286 163492 4338
rect 162988 4284 163492 4286
rect 163996 4340 164052 4350
rect 162988 4274 163044 4284
rect 163996 4246 164052 4284
rect 163324 4116 163380 4126
rect 162876 4060 163044 4116
rect 161756 4050 161812 4060
rect 161644 3826 161700 3836
rect 161532 3780 161588 3790
rect 161308 3778 161588 3780
rect 161308 3726 161534 3778
rect 161586 3726 161588 3778
rect 161308 3724 161588 3726
rect 161532 3714 161588 3724
rect 162316 3778 162372 3790
rect 162316 3726 162318 3778
rect 162370 3726 162372 3778
rect 162316 3668 162372 3726
rect 162316 3666 162708 3668
rect 162316 3614 162318 3666
rect 162370 3614 162708 3666
rect 162316 3612 162708 3614
rect 162316 3602 162372 3612
rect 162652 3554 162708 3612
rect 162652 3502 162654 3554
rect 162706 3502 162708 3554
rect 162652 3490 162708 3502
rect 161980 3444 162036 3482
rect 162988 3442 163044 4060
rect 162988 3390 162990 3442
rect 163042 3390 163044 3442
rect 161980 3332 162260 3388
rect 162988 3378 163044 3390
rect 163212 4114 163380 4116
rect 163212 4062 163326 4114
rect 163378 4062 163380 4114
rect 163212 4060 163380 4062
rect 160748 2706 160804 2716
rect 162204 800 162260 3332
rect 163212 2996 163268 4060
rect 163324 4050 163380 4060
rect 163324 3892 163380 3902
rect 163324 3442 163380 3836
rect 164332 3892 164388 5852
rect 164444 5906 164500 5918
rect 164444 5854 164446 5906
rect 164498 5854 164500 5906
rect 164444 5460 164500 5854
rect 164556 5572 164612 6188
rect 164556 5506 164612 5516
rect 164892 6130 164948 6636
rect 165116 6468 165172 6478
rect 165116 6374 165172 6412
rect 164892 6078 164894 6130
rect 164946 6078 164948 6130
rect 164444 5394 164500 5404
rect 164780 5348 164836 5358
rect 164780 5122 164836 5292
rect 164780 5070 164782 5122
rect 164834 5070 164836 5122
rect 164780 5058 164836 5070
rect 164892 5124 164948 6078
rect 165116 5908 165172 5918
rect 165116 5814 165172 5852
rect 165564 5908 165620 5918
rect 165564 5814 165620 5852
rect 165004 5794 165060 5806
rect 165004 5742 165006 5794
rect 165058 5742 165060 5794
rect 165004 5684 165060 5742
rect 165004 5618 165060 5628
rect 165676 5348 165732 5358
rect 165228 5236 165284 5246
rect 165228 5124 165284 5180
rect 164892 5122 165284 5124
rect 164892 5070 165230 5122
rect 165282 5070 165284 5122
rect 164892 5068 165284 5070
rect 165228 5058 165284 5068
rect 165676 5122 165732 5292
rect 165676 5070 165678 5122
rect 165730 5070 165732 5122
rect 165676 5058 165732 5070
rect 166124 5236 166180 5246
rect 166124 5122 166180 5180
rect 166124 5070 166126 5122
rect 166178 5070 166180 5122
rect 166124 5058 166180 5070
rect 166236 5124 166292 5134
rect 166236 5030 166292 5068
rect 164332 3826 164388 3836
rect 164444 4898 164500 4910
rect 164444 4846 164446 4898
rect 164498 4846 164500 4898
rect 163324 3390 163326 3442
rect 163378 3390 163380 3442
rect 163324 3378 163380 3390
rect 163660 3444 163716 3482
rect 163660 3378 163716 3388
rect 163212 2930 163268 2940
rect 164444 2884 164500 4846
rect 165340 4898 165396 4910
rect 165340 4846 165342 4898
rect 165394 4846 165396 4898
rect 165340 4452 165396 4846
rect 165452 4900 165508 4910
rect 166348 4900 166404 4910
rect 166908 4900 166964 4910
rect 165452 4898 165620 4900
rect 165452 4846 165454 4898
rect 165506 4846 165620 4898
rect 165452 4844 165620 4846
rect 165452 4834 165508 4844
rect 165340 4386 165396 4396
rect 165452 4340 165508 4350
rect 165004 3442 165060 3454
rect 165004 3390 165006 3442
rect 165058 3390 165060 3442
rect 165004 3388 165060 3390
rect 165452 3442 165508 4284
rect 165564 4228 165620 4844
rect 166348 4898 166964 4900
rect 166348 4846 166350 4898
rect 166402 4846 166910 4898
rect 166962 4846 166964 4898
rect 166348 4844 166964 4846
rect 166348 4834 166404 4844
rect 165676 4228 165732 4238
rect 165564 4172 165676 4228
rect 165676 4134 165732 4172
rect 166908 3668 166964 4844
rect 166908 3602 166964 3612
rect 165452 3390 165454 3442
rect 165506 3390 165508 3442
rect 164444 2818 164500 2828
rect 164892 3332 165396 3388
rect 165452 3378 165508 3390
rect 165676 3554 165732 3566
rect 165676 3502 165678 3554
rect 165730 3502 165732 3554
rect 164892 800 164948 3332
rect 165340 3220 165396 3332
rect 165676 3220 165732 3502
rect 165340 3164 165732 3220
rect 167580 3444 167636 3482
rect 167580 800 167636 3388
rect 167804 3330 167860 6748
rect 168140 3444 168196 3454
rect 168140 3350 168196 3388
rect 170268 3442 170324 3454
rect 170268 3390 170270 3442
rect 170322 3390 170324 3442
rect 167804 3278 167806 3330
rect 167858 3278 167860 3330
rect 167804 3266 167860 3278
rect 170268 3108 170324 3390
rect 170492 3330 170548 7308
rect 173436 6300 173700 6310
rect 173492 6244 173540 6300
rect 173596 6244 173644 6300
rect 173436 6234 173700 6244
rect 181244 5908 181300 5918
rect 178556 5012 178612 5022
rect 173436 4732 173700 4742
rect 173492 4676 173540 4732
rect 173596 4676 173644 4732
rect 173436 4666 173700 4676
rect 175868 3892 175924 3902
rect 173180 3780 173236 3790
rect 170492 3278 170494 3330
rect 170546 3278 170548 3330
rect 170492 3266 170548 3278
rect 170716 3554 170772 3566
rect 170716 3502 170718 3554
rect 170770 3502 170772 3554
rect 170716 3108 170772 3502
rect 172620 3444 172676 3454
rect 172956 3444 173012 3454
rect 172620 3442 172956 3444
rect 172620 3390 172622 3442
rect 172674 3390 172956 3442
rect 172620 3388 172956 3390
rect 172620 3378 172676 3388
rect 170268 3052 170772 3108
rect 170268 800 170324 3052
rect 172956 800 173012 3388
rect 173180 3442 173236 3724
rect 173180 3390 173182 3442
rect 173234 3390 173236 3442
rect 173180 3378 173236 3390
rect 173516 3444 173572 3454
rect 173516 3350 173572 3388
rect 175644 3442 175700 3454
rect 175644 3390 175646 3442
rect 175698 3390 175700 3442
rect 173436 3164 173700 3174
rect 173492 3108 173540 3164
rect 173596 3108 173644 3164
rect 173436 3098 173700 3108
rect 175644 3108 175700 3390
rect 175868 3330 175924 3836
rect 175868 3278 175870 3330
rect 175922 3278 175924 3330
rect 175868 3266 175924 3278
rect 176092 3554 176148 3566
rect 176092 3502 176094 3554
rect 176146 3502 176148 3554
rect 176092 3108 176148 3502
rect 175644 3052 176148 3108
rect 178332 3442 178388 3454
rect 178332 3390 178334 3442
rect 178386 3390 178388 3442
rect 178332 3108 178388 3390
rect 178556 3330 178612 4956
rect 178556 3278 178558 3330
rect 178610 3278 178612 3330
rect 178556 3266 178612 3278
rect 178780 3554 178836 3566
rect 178780 3502 178782 3554
rect 178834 3502 178836 3554
rect 178780 3108 178836 3502
rect 178332 3052 178836 3108
rect 181020 3444 181076 3454
rect 175644 800 175700 3052
rect 178332 800 178388 3052
rect 181020 800 181076 3388
rect 181244 3330 181300 5852
rect 181580 3444 181636 3454
rect 181580 3350 181636 3388
rect 181244 3278 181246 3330
rect 181298 3278 181300 3330
rect 181244 3266 181300 3278
rect 182252 2436 182308 45500
rect 184604 15988 184660 45614
rect 184604 15922 184660 15932
rect 187292 12964 187348 45724
rect 189196 45780 189252 45790
rect 189196 45686 189252 45724
rect 188796 44716 189060 44726
rect 188852 44660 188900 44716
rect 188956 44660 189004 44716
rect 188796 44650 189060 44660
rect 188796 43148 189060 43158
rect 188852 43092 188900 43148
rect 188956 43092 189004 43148
rect 188796 43082 189060 43092
rect 188796 41580 189060 41590
rect 188852 41524 188900 41580
rect 188956 41524 189004 41580
rect 188796 41514 189060 41524
rect 188796 40012 189060 40022
rect 188852 39956 188900 40012
rect 188956 39956 189004 40012
rect 188796 39946 189060 39956
rect 188796 38444 189060 38454
rect 188852 38388 188900 38444
rect 188956 38388 189004 38444
rect 188796 38378 189060 38388
rect 188796 36876 189060 36886
rect 188852 36820 188900 36876
rect 188956 36820 189004 36876
rect 188796 36810 189060 36820
rect 188796 35308 189060 35318
rect 188852 35252 188900 35308
rect 188956 35252 189004 35308
rect 188796 35242 189060 35252
rect 188796 33740 189060 33750
rect 188852 33684 188900 33740
rect 188956 33684 189004 33740
rect 188796 33674 189060 33684
rect 188796 32172 189060 32182
rect 188852 32116 188900 32172
rect 188956 32116 189004 32172
rect 188796 32106 189060 32116
rect 188796 30604 189060 30614
rect 188852 30548 188900 30604
rect 188956 30548 189004 30604
rect 188796 30538 189060 30548
rect 188796 29036 189060 29046
rect 188852 28980 188900 29036
rect 188956 28980 189004 29036
rect 188796 28970 189060 28980
rect 188796 27468 189060 27478
rect 188852 27412 188900 27468
rect 188956 27412 189004 27468
rect 188796 27402 189060 27412
rect 188796 25900 189060 25910
rect 188852 25844 188900 25900
rect 188956 25844 189004 25900
rect 188796 25834 189060 25844
rect 188796 24332 189060 24342
rect 188852 24276 188900 24332
rect 188956 24276 189004 24332
rect 188796 24266 189060 24276
rect 188796 22764 189060 22774
rect 188852 22708 188900 22764
rect 188956 22708 189004 22764
rect 188796 22698 189060 22708
rect 188796 21196 189060 21206
rect 188852 21140 188900 21196
rect 188956 21140 189004 21196
rect 188796 21130 189060 21140
rect 188796 19628 189060 19638
rect 188852 19572 188900 19628
rect 188956 19572 189004 19628
rect 188796 19562 189060 19572
rect 188796 18060 189060 18070
rect 188852 18004 188900 18060
rect 188956 18004 189004 18060
rect 188796 17994 189060 18004
rect 188796 16492 189060 16502
rect 188852 16436 188900 16492
rect 188956 16436 189004 16492
rect 188796 16426 189060 16436
rect 188796 14924 189060 14934
rect 188852 14868 188900 14924
rect 188956 14868 189004 14924
rect 188796 14858 189060 14868
rect 188796 13356 189060 13366
rect 188852 13300 188900 13356
rect 188956 13300 189004 13356
rect 188796 13290 189060 13300
rect 187292 12898 187348 12908
rect 193116 12852 193172 45950
rect 196476 46004 196532 49200
rect 200508 46004 200564 49200
rect 204540 46004 204596 49200
rect 205212 46004 205268 46014
rect 196476 46002 196756 46004
rect 196476 45950 196478 46002
rect 196530 45950 196756 46002
rect 196476 45948 196756 45950
rect 196476 45910 196532 45948
rect 196700 45890 196756 45948
rect 200508 46002 200788 46004
rect 200508 45950 200510 46002
rect 200562 45950 200788 46002
rect 200508 45948 200788 45950
rect 200508 45938 200564 45948
rect 196700 45838 196702 45890
rect 196754 45838 196756 45890
rect 196700 45826 196756 45838
rect 200732 45890 200788 45948
rect 204540 46002 204820 46004
rect 204540 45950 204542 46002
rect 204594 45950 204820 46002
rect 204540 45948 204820 45950
rect 204540 45938 204596 45948
rect 200732 45838 200734 45890
rect 200786 45838 200788 45890
rect 200732 45826 200788 45838
rect 204764 45890 204820 45948
rect 205212 45910 205268 45948
rect 205772 46004 205828 46014
rect 204764 45838 204766 45890
rect 204818 45838 204820 45890
rect 204764 45826 204820 45838
rect 197260 45778 197316 45790
rect 197260 45726 197262 45778
rect 197314 45726 197316 45778
rect 197260 17668 197316 45726
rect 201292 45780 201348 45790
rect 201292 45686 201348 45724
rect 204156 45500 204420 45510
rect 204212 45444 204260 45500
rect 204316 45444 204364 45500
rect 204156 45434 204420 45444
rect 204156 43932 204420 43942
rect 204212 43876 204260 43932
rect 204316 43876 204364 43932
rect 204156 43866 204420 43876
rect 204156 42364 204420 42374
rect 204212 42308 204260 42364
rect 204316 42308 204364 42364
rect 204156 42298 204420 42308
rect 204156 40796 204420 40806
rect 204212 40740 204260 40796
rect 204316 40740 204364 40796
rect 204156 40730 204420 40740
rect 204156 39228 204420 39238
rect 204212 39172 204260 39228
rect 204316 39172 204364 39228
rect 204156 39162 204420 39172
rect 204156 37660 204420 37670
rect 204212 37604 204260 37660
rect 204316 37604 204364 37660
rect 204156 37594 204420 37604
rect 204156 36092 204420 36102
rect 204212 36036 204260 36092
rect 204316 36036 204364 36092
rect 204156 36026 204420 36036
rect 204156 34524 204420 34534
rect 204212 34468 204260 34524
rect 204316 34468 204364 34524
rect 204156 34458 204420 34468
rect 204156 32956 204420 32966
rect 204212 32900 204260 32956
rect 204316 32900 204364 32956
rect 204156 32890 204420 32900
rect 204156 31388 204420 31398
rect 204212 31332 204260 31388
rect 204316 31332 204364 31388
rect 204156 31322 204420 31332
rect 204156 29820 204420 29830
rect 204212 29764 204260 29820
rect 204316 29764 204364 29820
rect 204156 29754 204420 29764
rect 204156 28252 204420 28262
rect 204212 28196 204260 28252
rect 204316 28196 204364 28252
rect 204156 28186 204420 28196
rect 204156 26684 204420 26694
rect 204212 26628 204260 26684
rect 204316 26628 204364 26684
rect 204156 26618 204420 26628
rect 204156 25116 204420 25126
rect 204212 25060 204260 25116
rect 204316 25060 204364 25116
rect 204156 25050 204420 25060
rect 204156 23548 204420 23558
rect 204212 23492 204260 23548
rect 204316 23492 204364 23548
rect 204156 23482 204420 23492
rect 204156 21980 204420 21990
rect 204212 21924 204260 21980
rect 204316 21924 204364 21980
rect 204156 21914 204420 21924
rect 204156 20412 204420 20422
rect 204212 20356 204260 20412
rect 204316 20356 204364 20412
rect 204156 20346 204420 20356
rect 204156 18844 204420 18854
rect 204212 18788 204260 18844
rect 204316 18788 204364 18844
rect 204156 18778 204420 18788
rect 197260 17602 197316 17612
rect 204156 17276 204420 17286
rect 204212 17220 204260 17276
rect 204316 17220 204364 17276
rect 204156 17210 204420 17220
rect 204156 15708 204420 15718
rect 204212 15652 204260 15708
rect 204316 15652 204364 15708
rect 204156 15642 204420 15652
rect 204156 14140 204420 14150
rect 204212 14084 204260 14140
rect 204316 14084 204364 14140
rect 204156 14074 204420 14084
rect 193116 12786 193172 12796
rect 204156 12572 204420 12582
rect 204212 12516 204260 12572
rect 204316 12516 204364 12572
rect 204156 12506 204420 12516
rect 188796 11788 189060 11798
rect 188852 11732 188900 11788
rect 188956 11732 189004 11788
rect 188796 11722 189060 11732
rect 204156 11004 204420 11014
rect 204212 10948 204260 11004
rect 204316 10948 204364 11004
rect 204156 10938 204420 10948
rect 188796 10220 189060 10230
rect 188852 10164 188900 10220
rect 188956 10164 189004 10220
rect 188796 10154 189060 10164
rect 204156 9436 204420 9446
rect 204212 9380 204260 9436
rect 204316 9380 204364 9436
rect 204156 9370 204420 9380
rect 188796 8652 189060 8662
rect 188852 8596 188900 8652
rect 188956 8596 189004 8652
rect 188796 8586 189060 8596
rect 204156 7868 204420 7878
rect 204212 7812 204260 7868
rect 204316 7812 204364 7868
rect 204156 7802 204420 7812
rect 205772 7700 205828 45948
rect 208572 46004 208628 49200
rect 212604 46004 212660 49200
rect 216636 46004 216692 49200
rect 217532 46004 217588 46014
rect 208572 46002 208852 46004
rect 208572 45950 208574 46002
rect 208626 45950 208852 46002
rect 208572 45948 208852 45950
rect 208572 45938 208628 45948
rect 208796 45890 208852 45948
rect 212604 46002 212884 46004
rect 212604 45950 212606 46002
rect 212658 45950 212884 46002
rect 212604 45948 212884 45950
rect 212604 45938 212660 45948
rect 208796 45838 208798 45890
rect 208850 45838 208852 45890
rect 208796 45826 208852 45838
rect 212828 45890 212884 45948
rect 216636 46002 216916 46004
rect 216636 45950 216638 46002
rect 216690 45950 216916 46002
rect 216636 45948 216916 45950
rect 216636 45938 216692 45948
rect 212828 45838 212830 45890
rect 212882 45838 212884 45890
rect 212828 45826 212884 45838
rect 216860 45890 216916 45948
rect 217532 45910 217588 45948
rect 216860 45838 216862 45890
rect 216914 45838 216916 45890
rect 216860 45826 216916 45838
rect 209356 45778 209412 45790
rect 209356 45726 209358 45778
rect 209410 45726 209412 45778
rect 209356 14308 209412 45726
rect 209356 14242 209412 14252
rect 213948 45778 214004 45790
rect 213948 45726 213950 45778
rect 214002 45726 214004 45778
rect 213948 12740 214004 45726
rect 213948 12674 214004 12684
rect 205772 7634 205828 7644
rect 188796 7084 189060 7094
rect 188852 7028 188900 7084
rect 188956 7028 189004 7084
rect 188796 7018 189060 7028
rect 213948 6916 214004 6926
rect 204156 6300 204420 6310
rect 204212 6244 204260 6300
rect 204316 6244 204364 6300
rect 204156 6234 204420 6244
rect 189308 6132 189364 6142
rect 188796 5516 189060 5526
rect 188852 5460 188900 5516
rect 188956 5460 189004 5516
rect 188796 5450 189060 5460
rect 184492 4228 184548 4238
rect 182252 2370 182308 2380
rect 184044 3442 184100 3454
rect 184044 3390 184046 3442
rect 184098 3390 184100 3442
rect 184044 3108 184100 3390
rect 184492 3330 184548 4172
rect 188796 3948 189060 3958
rect 188852 3892 188900 3948
rect 188956 3892 189004 3948
rect 188796 3882 189060 3892
rect 186620 3780 186676 3790
rect 184492 3278 184494 3330
rect 184546 3278 184548 3330
rect 184492 3266 184548 3278
rect 184716 3554 184772 3566
rect 184716 3502 184718 3554
rect 184770 3502 184772 3554
rect 184716 3108 184772 3502
rect 184044 3052 184772 3108
rect 186396 3444 186452 3454
rect 184044 2324 184100 3052
rect 183708 2268 184100 2324
rect 183708 800 183764 2268
rect 186396 800 186452 3388
rect 186620 3330 186676 3724
rect 186844 3554 186900 3566
rect 186844 3502 186846 3554
rect 186898 3502 186900 3554
rect 186844 3444 186900 3502
rect 186844 3378 186900 3388
rect 189084 3442 189140 3454
rect 189084 3390 189086 3442
rect 189138 3390 189140 3442
rect 186620 3278 186622 3330
rect 186674 3278 186676 3330
rect 186620 3266 186676 3278
rect 189084 3108 189140 3390
rect 189308 3330 189364 6076
rect 192108 6020 192164 6030
rect 189308 3278 189310 3330
rect 189362 3278 189364 3330
rect 189308 3266 189364 3278
rect 189532 3554 189588 3566
rect 189532 3502 189534 3554
rect 189586 3502 189588 3554
rect 189532 3108 189588 3502
rect 191660 3444 191716 3454
rect 191660 3442 191828 3444
rect 191660 3390 191662 3442
rect 191714 3390 191828 3442
rect 191660 3388 191828 3390
rect 191660 3378 191716 3388
rect 189084 3052 189588 3108
rect 191772 3108 191828 3388
rect 192108 3330 192164 5964
rect 194684 5684 194740 5694
rect 192108 3278 192110 3330
rect 192162 3278 192164 3330
rect 192108 3266 192164 3278
rect 192332 3554 192388 3566
rect 192332 3502 192334 3554
rect 192386 3502 192388 3554
rect 192332 3108 192388 3502
rect 191772 3052 192388 3108
rect 194460 3444 194516 3454
rect 189084 800 189140 3052
rect 191772 800 191828 3052
rect 194460 800 194516 3388
rect 194684 3330 194740 5628
rect 204156 4732 204420 4742
rect 204212 4676 204260 4732
rect 204316 4676 204364 4732
rect 204156 4666 204420 4676
rect 211596 3668 211652 3678
rect 211596 3574 211652 3612
rect 213948 3666 214004 6860
rect 213948 3614 213950 3666
rect 214002 3614 214004 3666
rect 213948 3602 214004 3614
rect 216636 4564 216692 4574
rect 216636 3666 216692 4508
rect 216636 3614 216638 3666
rect 216690 3614 216692 3666
rect 216636 3602 216692 3614
rect 197932 3554 197988 3566
rect 197932 3502 197934 3554
rect 197986 3502 197988 3554
rect 195020 3444 195076 3454
rect 195020 3350 195076 3388
rect 197148 3444 197204 3454
rect 197372 3444 197428 3454
rect 197148 3442 197428 3444
rect 197148 3390 197150 3442
rect 197202 3390 197374 3442
rect 197426 3390 197428 3442
rect 197148 3388 197428 3390
rect 194684 3278 194686 3330
rect 194738 3278 194740 3330
rect 194684 3266 194740 3278
rect 197148 800 197204 3388
rect 197372 3378 197428 3388
rect 197932 2212 197988 3502
rect 205996 3554 206052 3566
rect 205996 3502 205998 3554
rect 206050 3502 206052 3554
rect 199276 3444 199332 3454
rect 200060 3444 200116 3454
rect 199276 3442 200116 3444
rect 199276 3390 199278 3442
rect 199330 3390 200062 3442
rect 200114 3390 200116 3442
rect 199276 3388 200116 3390
rect 199276 3378 199332 3388
rect 197932 2146 197988 2156
rect 199836 800 199892 3388
rect 200060 3378 200116 3388
rect 200620 3442 200676 3454
rect 200620 3390 200622 3442
rect 200674 3390 200676 3442
rect 200620 1428 200676 3390
rect 203084 3444 203140 3454
rect 203532 3444 203588 3454
rect 204092 3444 204148 3454
rect 203084 3442 203588 3444
rect 203084 3390 203086 3442
rect 203138 3390 203534 3442
rect 203586 3390 203588 3442
rect 203084 3388 203588 3390
rect 203084 2212 203140 3388
rect 203532 3378 203588 3388
rect 203980 3442 204148 3444
rect 203980 3390 204094 3442
rect 204146 3390 204148 3442
rect 203980 3388 204148 3390
rect 200620 1362 200676 1372
rect 202524 2156 203140 2212
rect 202524 800 202580 2156
rect 203980 1652 204036 3388
rect 204092 3378 204148 3388
rect 205212 3444 205268 3454
rect 205436 3444 205492 3454
rect 205212 3442 205492 3444
rect 205212 3390 205214 3442
rect 205266 3390 205438 3442
rect 205490 3390 205492 3442
rect 205212 3388 205492 3390
rect 204156 3164 204420 3174
rect 204212 3108 204260 3164
rect 204316 3108 204364 3164
rect 204156 3098 204420 3108
rect 203980 1586 204036 1596
rect 205212 800 205268 3388
rect 205436 3378 205492 3388
rect 205996 3332 206052 3502
rect 205996 3266 206052 3276
rect 207900 3444 207956 3454
rect 208124 3444 208180 3454
rect 207900 3442 208180 3444
rect 207900 3390 207902 3442
rect 207954 3390 208126 3442
rect 208178 3390 208180 3442
rect 207900 3388 208180 3390
rect 207900 800 207956 3388
rect 208124 3378 208180 3388
rect 208684 3442 208740 3454
rect 210700 3444 210756 3454
rect 211148 3444 211204 3454
rect 208684 3390 208686 3442
rect 208738 3390 208740 3442
rect 208684 1540 208740 3390
rect 208684 1474 208740 1484
rect 210588 3442 211204 3444
rect 210588 3390 210702 3442
rect 210754 3390 211150 3442
rect 211202 3390 211204 3442
rect 210588 3388 211204 3390
rect 210588 800 210644 3388
rect 210700 3378 210756 3388
rect 211148 3378 211204 3388
rect 213276 3444 213332 3454
rect 213500 3444 213556 3454
rect 213276 3442 213556 3444
rect 213276 3390 213278 3442
rect 213330 3390 213502 3442
rect 213554 3390 213556 3442
rect 213276 3388 213556 3390
rect 213276 800 213332 3388
rect 213500 3378 213556 3388
rect 215964 3444 216020 3454
rect 216188 3444 216244 3454
rect 215964 3442 216244 3444
rect 215964 3390 215966 3442
rect 216018 3390 216190 3442
rect 216242 3390 216244 3442
rect 215964 3388 216244 3390
rect 215964 800 216020 3388
rect 216188 3378 216244 3388
rect 3584 0 3696 800
rect 6272 0 6384 800
rect 8960 0 9072 800
rect 11648 0 11760 800
rect 14336 0 14448 800
rect 17024 0 17136 800
rect 19712 0 19824 800
rect 22400 0 22512 800
rect 25088 0 25200 800
rect 27776 0 27888 800
rect 30464 0 30576 800
rect 33152 0 33264 800
rect 35840 0 35952 800
rect 38528 0 38640 800
rect 41216 0 41328 800
rect 43904 0 44016 800
rect 46592 0 46704 800
rect 49280 0 49392 800
rect 51968 0 52080 800
rect 54656 0 54768 800
rect 57344 0 57456 800
rect 60032 0 60144 800
rect 62720 0 62832 800
rect 65408 0 65520 800
rect 68096 0 68208 800
rect 70784 0 70896 800
rect 73472 0 73584 800
rect 76160 0 76272 800
rect 78848 0 78960 800
rect 81536 0 81648 800
rect 84224 0 84336 800
rect 86912 0 87024 800
rect 89600 0 89712 800
rect 92288 0 92400 800
rect 94976 0 95088 800
rect 97664 0 97776 800
rect 100352 0 100464 800
rect 103040 0 103152 800
rect 105728 0 105840 800
rect 108416 0 108528 800
rect 111104 0 111216 800
rect 113792 0 113904 800
rect 116480 0 116592 800
rect 119168 0 119280 800
rect 121856 0 121968 800
rect 124544 0 124656 800
rect 127232 0 127344 800
rect 129920 0 130032 800
rect 132608 0 132720 800
rect 135296 0 135408 800
rect 137984 0 138096 800
rect 140672 0 140784 800
rect 143360 0 143472 800
rect 146048 0 146160 800
rect 148736 0 148848 800
rect 151424 0 151536 800
rect 154112 0 154224 800
rect 156800 0 156912 800
rect 159488 0 159600 800
rect 162176 0 162288 800
rect 164864 0 164976 800
rect 167552 0 167664 800
rect 170240 0 170352 800
rect 172928 0 173040 800
rect 175616 0 175728 800
rect 178304 0 178416 800
rect 180992 0 181104 800
rect 183680 0 183792 800
rect 186368 0 186480 800
rect 189056 0 189168 800
rect 191744 0 191856 800
rect 194432 0 194544 800
rect 197120 0 197232 800
rect 199808 0 199920 800
rect 202496 0 202608 800
rect 205184 0 205296 800
rect 207872 0 207984 800
rect 210560 0 210672 800
rect 213248 0 213360 800
rect 215936 0 216048 800
<< via2 >>
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 2940 37100 2996 37156
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 5964 5180 6020 5236
rect 6412 5234 6468 5236
rect 6412 5182 6414 5234
rect 6414 5182 6466 5234
rect 6466 5182 6468 5234
rect 6412 5180 6468 5182
rect 12348 45052 12404 45108
rect 19852 45890 19908 45892
rect 19852 45838 19854 45890
rect 19854 45838 19906 45890
rect 19906 45838 19908 45890
rect 19852 45836 19908 45838
rect 22652 45836 22708 45892
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 31612 46002 31668 46004
rect 31612 45950 31614 46002
rect 31614 45950 31666 46002
rect 31666 45950 31668 46002
rect 31612 45948 31668 45950
rect 32172 45948 32228 46004
rect 23884 26012 23940 26068
rect 36540 45890 36596 45892
rect 36540 45838 36542 45890
rect 36542 45838 36594 45890
rect 36594 45838 36596 45890
rect 36540 45836 36596 45838
rect 37772 45836 37828 45892
rect 32732 45388 32788 45444
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 37772 15932 37828 15988
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 28924 12684 28980 12740
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 65916 46282 65972 46284
rect 65916 46230 65918 46282
rect 65918 46230 65970 46282
rect 65970 46230 65972 46282
rect 65916 46228 65972 46230
rect 66020 46282 66076 46284
rect 66020 46230 66022 46282
rect 66022 46230 66074 46282
rect 66074 46230 66076 46282
rect 66020 46228 66076 46230
rect 66124 46282 66180 46284
rect 66124 46230 66126 46282
rect 66126 46230 66178 46282
rect 66178 46230 66180 46282
rect 66124 46228 66180 46230
rect 44156 45890 44212 45892
rect 44156 45838 44158 45890
rect 44158 45838 44210 45890
rect 44210 45838 44212 45890
rect 44156 45836 44212 45838
rect 47852 45836 47908 45892
rect 42812 45388 42868 45444
rect 54124 45890 54180 45892
rect 54124 45838 54126 45890
rect 54126 45838 54178 45890
rect 54178 45838 54180 45890
rect 54124 45836 54180 45838
rect 55132 45890 55188 45892
rect 55132 45838 55134 45890
rect 55134 45838 55186 45890
rect 55186 45838 55188 45890
rect 55132 45836 55188 45838
rect 58044 45836 58100 45892
rect 50092 45612 50148 45668
rect 50540 45666 50596 45668
rect 50540 45614 50542 45666
rect 50542 45614 50594 45666
rect 50594 45614 50596 45666
rect 50540 45612 50596 45614
rect 52892 45612 52948 45668
rect 50556 45498 50612 45500
rect 50556 45446 50558 45498
rect 50558 45446 50610 45498
rect 50610 45446 50612 45498
rect 50556 45444 50612 45446
rect 50660 45498 50716 45500
rect 50660 45446 50662 45498
rect 50662 45446 50714 45498
rect 50714 45446 50716 45498
rect 50660 45444 50716 45446
rect 50764 45498 50820 45500
rect 50764 45446 50766 45498
rect 50766 45446 50818 45498
rect 50818 45446 50820 45498
rect 50764 45444 50820 45446
rect 50556 43930 50612 43932
rect 50556 43878 50558 43930
rect 50558 43878 50610 43930
rect 50610 43878 50612 43930
rect 50556 43876 50612 43878
rect 50660 43930 50716 43932
rect 50660 43878 50662 43930
rect 50662 43878 50714 43930
rect 50714 43878 50716 43930
rect 50660 43876 50716 43878
rect 50764 43930 50820 43932
rect 50764 43878 50766 43930
rect 50766 43878 50818 43930
rect 50818 43878 50820 43930
rect 50764 43876 50820 43878
rect 50556 42362 50612 42364
rect 50556 42310 50558 42362
rect 50558 42310 50610 42362
rect 50610 42310 50612 42362
rect 50556 42308 50612 42310
rect 50660 42362 50716 42364
rect 50660 42310 50662 42362
rect 50662 42310 50714 42362
rect 50714 42310 50716 42362
rect 50660 42308 50716 42310
rect 50764 42362 50820 42364
rect 50764 42310 50766 42362
rect 50766 42310 50818 42362
rect 50818 42310 50820 42362
rect 50764 42308 50820 42310
rect 50556 40794 50612 40796
rect 50556 40742 50558 40794
rect 50558 40742 50610 40794
rect 50610 40742 50612 40794
rect 50556 40740 50612 40742
rect 50660 40794 50716 40796
rect 50660 40742 50662 40794
rect 50662 40742 50714 40794
rect 50714 40742 50716 40794
rect 50660 40740 50716 40742
rect 50764 40794 50820 40796
rect 50764 40742 50766 40794
rect 50766 40742 50818 40794
rect 50818 40742 50820 40794
rect 50764 40740 50820 40742
rect 50556 39226 50612 39228
rect 50556 39174 50558 39226
rect 50558 39174 50610 39226
rect 50610 39174 50612 39226
rect 50556 39172 50612 39174
rect 50660 39226 50716 39228
rect 50660 39174 50662 39226
rect 50662 39174 50714 39226
rect 50714 39174 50716 39226
rect 50660 39172 50716 39174
rect 50764 39226 50820 39228
rect 50764 39174 50766 39226
rect 50766 39174 50818 39226
rect 50818 39174 50820 39226
rect 50764 39172 50820 39174
rect 50556 37658 50612 37660
rect 50556 37606 50558 37658
rect 50558 37606 50610 37658
rect 50610 37606 50612 37658
rect 50556 37604 50612 37606
rect 50660 37658 50716 37660
rect 50660 37606 50662 37658
rect 50662 37606 50714 37658
rect 50714 37606 50716 37658
rect 50660 37604 50716 37606
rect 50764 37658 50820 37660
rect 50764 37606 50766 37658
rect 50766 37606 50818 37658
rect 50818 37606 50820 37658
rect 50764 37604 50820 37606
rect 50556 36090 50612 36092
rect 50556 36038 50558 36090
rect 50558 36038 50610 36090
rect 50610 36038 50612 36090
rect 50556 36036 50612 36038
rect 50660 36090 50716 36092
rect 50660 36038 50662 36090
rect 50662 36038 50714 36090
rect 50714 36038 50716 36090
rect 50660 36036 50716 36038
rect 50764 36090 50820 36092
rect 50764 36038 50766 36090
rect 50766 36038 50818 36090
rect 50818 36038 50820 36090
rect 50764 36036 50820 36038
rect 50556 34522 50612 34524
rect 50556 34470 50558 34522
rect 50558 34470 50610 34522
rect 50610 34470 50612 34522
rect 50556 34468 50612 34470
rect 50660 34522 50716 34524
rect 50660 34470 50662 34522
rect 50662 34470 50714 34522
rect 50714 34470 50716 34522
rect 50660 34468 50716 34470
rect 50764 34522 50820 34524
rect 50764 34470 50766 34522
rect 50766 34470 50818 34522
rect 50818 34470 50820 34522
rect 50764 34468 50820 34470
rect 50556 32954 50612 32956
rect 50556 32902 50558 32954
rect 50558 32902 50610 32954
rect 50610 32902 50612 32954
rect 50556 32900 50612 32902
rect 50660 32954 50716 32956
rect 50660 32902 50662 32954
rect 50662 32902 50714 32954
rect 50714 32902 50716 32954
rect 50660 32900 50716 32902
rect 50764 32954 50820 32956
rect 50764 32902 50766 32954
rect 50766 32902 50818 32954
rect 50818 32902 50820 32954
rect 50764 32900 50820 32902
rect 50556 31386 50612 31388
rect 50556 31334 50558 31386
rect 50558 31334 50610 31386
rect 50610 31334 50612 31386
rect 50556 31332 50612 31334
rect 50660 31386 50716 31388
rect 50660 31334 50662 31386
rect 50662 31334 50714 31386
rect 50714 31334 50716 31386
rect 50660 31332 50716 31334
rect 50764 31386 50820 31388
rect 50764 31334 50766 31386
rect 50766 31334 50818 31386
rect 50818 31334 50820 31386
rect 50764 31332 50820 31334
rect 50556 29818 50612 29820
rect 50556 29766 50558 29818
rect 50558 29766 50610 29818
rect 50610 29766 50612 29818
rect 50556 29764 50612 29766
rect 50660 29818 50716 29820
rect 50660 29766 50662 29818
rect 50662 29766 50714 29818
rect 50714 29766 50716 29818
rect 50660 29764 50716 29766
rect 50764 29818 50820 29820
rect 50764 29766 50766 29818
rect 50766 29766 50818 29818
rect 50818 29766 50820 29818
rect 50764 29764 50820 29766
rect 50556 28250 50612 28252
rect 50556 28198 50558 28250
rect 50558 28198 50610 28250
rect 50610 28198 50612 28250
rect 50556 28196 50612 28198
rect 50660 28250 50716 28252
rect 50660 28198 50662 28250
rect 50662 28198 50714 28250
rect 50714 28198 50716 28250
rect 50660 28196 50716 28198
rect 50764 28250 50820 28252
rect 50764 28198 50766 28250
rect 50766 28198 50818 28250
rect 50818 28198 50820 28250
rect 50764 28196 50820 28198
rect 50556 26682 50612 26684
rect 50556 26630 50558 26682
rect 50558 26630 50610 26682
rect 50610 26630 50612 26682
rect 50556 26628 50612 26630
rect 50660 26682 50716 26684
rect 50660 26630 50662 26682
rect 50662 26630 50714 26682
rect 50714 26630 50716 26682
rect 50660 26628 50716 26630
rect 50764 26682 50820 26684
rect 50764 26630 50766 26682
rect 50766 26630 50818 26682
rect 50818 26630 50820 26682
rect 50764 26628 50820 26630
rect 50556 25114 50612 25116
rect 50556 25062 50558 25114
rect 50558 25062 50610 25114
rect 50610 25062 50612 25114
rect 50556 25060 50612 25062
rect 50660 25114 50716 25116
rect 50660 25062 50662 25114
rect 50662 25062 50714 25114
rect 50714 25062 50716 25114
rect 50660 25060 50716 25062
rect 50764 25114 50820 25116
rect 50764 25062 50766 25114
rect 50766 25062 50818 25114
rect 50818 25062 50820 25114
rect 50764 25060 50820 25062
rect 50556 23546 50612 23548
rect 50556 23494 50558 23546
rect 50558 23494 50610 23546
rect 50610 23494 50612 23546
rect 50556 23492 50612 23494
rect 50660 23546 50716 23548
rect 50660 23494 50662 23546
rect 50662 23494 50714 23546
rect 50714 23494 50716 23546
rect 50660 23492 50716 23494
rect 50764 23546 50820 23548
rect 50764 23494 50766 23546
rect 50766 23494 50818 23546
rect 50818 23494 50820 23546
rect 50764 23492 50820 23494
rect 50556 21978 50612 21980
rect 50556 21926 50558 21978
rect 50558 21926 50610 21978
rect 50610 21926 50612 21978
rect 50556 21924 50612 21926
rect 50660 21978 50716 21980
rect 50660 21926 50662 21978
rect 50662 21926 50714 21978
rect 50714 21926 50716 21978
rect 50660 21924 50716 21926
rect 50764 21978 50820 21980
rect 50764 21926 50766 21978
rect 50766 21926 50818 21978
rect 50818 21926 50820 21978
rect 50764 21924 50820 21926
rect 50556 20410 50612 20412
rect 50556 20358 50558 20410
rect 50558 20358 50610 20410
rect 50610 20358 50612 20410
rect 50556 20356 50612 20358
rect 50660 20410 50716 20412
rect 50660 20358 50662 20410
rect 50662 20358 50714 20410
rect 50714 20358 50716 20410
rect 50660 20356 50716 20358
rect 50764 20410 50820 20412
rect 50764 20358 50766 20410
rect 50766 20358 50818 20410
rect 50818 20358 50820 20410
rect 50764 20356 50820 20358
rect 47852 19292 47908 19348
rect 50556 18842 50612 18844
rect 50556 18790 50558 18842
rect 50558 18790 50610 18842
rect 50610 18790 50612 18842
rect 50556 18788 50612 18790
rect 50660 18842 50716 18844
rect 50660 18790 50662 18842
rect 50662 18790 50714 18842
rect 50714 18790 50716 18842
rect 50660 18788 50716 18790
rect 50764 18842 50820 18844
rect 50764 18790 50766 18842
rect 50766 18790 50818 18842
rect 50818 18790 50820 18842
rect 50764 18788 50820 18790
rect 50556 17274 50612 17276
rect 50556 17222 50558 17274
rect 50558 17222 50610 17274
rect 50610 17222 50612 17274
rect 50556 17220 50612 17222
rect 50660 17274 50716 17276
rect 50660 17222 50662 17274
rect 50662 17222 50714 17274
rect 50714 17222 50716 17274
rect 50660 17220 50716 17222
rect 50764 17274 50820 17276
rect 50764 17222 50766 17274
rect 50766 17222 50818 17274
rect 50818 17222 50820 17274
rect 50764 17220 50820 17222
rect 50556 15706 50612 15708
rect 50556 15654 50558 15706
rect 50558 15654 50610 15706
rect 50610 15654 50612 15706
rect 50556 15652 50612 15654
rect 50660 15706 50716 15708
rect 50660 15654 50662 15706
rect 50662 15654 50714 15706
rect 50714 15654 50716 15706
rect 50660 15652 50716 15654
rect 50764 15706 50820 15708
rect 50764 15654 50766 15706
rect 50766 15654 50818 15706
rect 50818 15654 50820 15706
rect 50764 15652 50820 15654
rect 42812 14252 42868 14308
rect 50556 14138 50612 14140
rect 50556 14086 50558 14138
rect 50558 14086 50610 14138
rect 50610 14086 50612 14138
rect 50556 14084 50612 14086
rect 50660 14138 50716 14140
rect 50660 14086 50662 14138
rect 50662 14086 50714 14138
rect 50714 14086 50716 14138
rect 50660 14084 50716 14086
rect 50764 14138 50820 14140
rect 50764 14086 50766 14138
rect 50766 14086 50818 14138
rect 50818 14086 50820 14138
rect 50764 14084 50820 14086
rect 50556 12570 50612 12572
rect 50556 12518 50558 12570
rect 50558 12518 50610 12570
rect 50610 12518 50612 12570
rect 50556 12516 50612 12518
rect 50660 12570 50716 12572
rect 50660 12518 50662 12570
rect 50662 12518 50714 12570
rect 50714 12518 50716 12570
rect 50660 12516 50716 12518
rect 50764 12570 50820 12572
rect 50764 12518 50766 12570
rect 50766 12518 50818 12570
rect 50818 12518 50820 12570
rect 50764 12516 50820 12518
rect 40236 11228 40292 11284
rect 52892 11116 52948 11172
rect 55132 26012 55188 26068
rect 50556 11002 50612 11004
rect 50556 10950 50558 11002
rect 50558 10950 50610 11002
rect 50610 10950 50612 11002
rect 50556 10948 50612 10950
rect 50660 11002 50716 11004
rect 50660 10950 50662 11002
rect 50662 10950 50714 11002
rect 50714 10950 50716 11002
rect 50660 10948 50716 10950
rect 50764 11002 50820 11004
rect 50764 10950 50766 11002
rect 50766 10950 50818 11002
rect 50818 10950 50820 11002
rect 50764 10948 50820 10950
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 50556 9434 50612 9436
rect 50556 9382 50558 9434
rect 50558 9382 50610 9434
rect 50610 9382 50612 9434
rect 50556 9380 50612 9382
rect 50660 9434 50716 9436
rect 50660 9382 50662 9434
rect 50662 9382 50714 9434
rect 50714 9382 50716 9434
rect 50660 9380 50716 9382
rect 50764 9434 50820 9436
rect 50764 9382 50766 9434
rect 50766 9382 50818 9434
rect 50818 9382 50820 9434
rect 50764 9380 50820 9382
rect 22652 9212 22708 9268
rect 52108 9212 52164 9268
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 50556 7866 50612 7868
rect 50556 7814 50558 7866
rect 50558 7814 50610 7866
rect 50610 7814 50612 7866
rect 50556 7812 50612 7814
rect 50660 7866 50716 7868
rect 50660 7814 50662 7866
rect 50662 7814 50714 7866
rect 50714 7814 50716 7866
rect 50660 7812 50716 7814
rect 50764 7866 50820 7868
rect 50764 7814 50766 7866
rect 50766 7814 50818 7866
rect 50818 7814 50820 7866
rect 50764 7812 50820 7814
rect 15820 7532 15876 7588
rect 49756 7532 49812 7588
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 33180 6860 33236 6916
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 7196 5180 7252 5236
rect 31500 5740 31556 5796
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 27804 3612 27860 3668
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 28588 3666 28644 3668
rect 28588 3614 28590 3666
rect 28590 3614 28642 3666
rect 28642 3614 28644 3666
rect 28588 3612 28644 3614
rect 39228 6748 39284 6804
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 35644 4562 35700 4564
rect 35644 4510 35646 4562
rect 35646 4510 35698 4562
rect 35698 4510 35700 4562
rect 35644 4508 35700 4510
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 44492 5964 44548 6020
rect 50556 6298 50612 6300
rect 50556 6246 50558 6298
rect 50558 6246 50610 6298
rect 50610 6246 50612 6298
rect 50556 6244 50612 6246
rect 50660 6298 50716 6300
rect 50660 6246 50662 6298
rect 50662 6246 50714 6298
rect 50714 6246 50716 6298
rect 50660 6244 50716 6246
rect 50764 6298 50820 6300
rect 50764 6246 50766 6298
rect 50766 6246 50818 6298
rect 50818 6246 50820 6298
rect 50764 6244 50820 6246
rect 57820 12684 57876 12740
rect 57036 5852 57092 5908
rect 46956 4844 47012 4900
rect 38556 3388 38612 3444
rect 40572 3442 40628 3444
rect 40572 3390 40574 3442
rect 40574 3390 40626 3442
rect 40626 3390 40628 3442
rect 40572 3388 40628 3390
rect 42364 3612 42420 3668
rect 42924 3666 42980 3668
rect 42924 3614 42926 3666
rect 42926 3614 42978 3666
rect 42978 3614 42980 3666
rect 42924 3612 42980 3614
rect 49980 4172 50036 4228
rect 46620 3388 46676 3444
rect 47628 3388 47684 3444
rect 50556 4730 50612 4732
rect 50556 4678 50558 4730
rect 50558 4678 50610 4730
rect 50610 4678 50612 4730
rect 50556 4676 50612 4678
rect 50660 4730 50716 4732
rect 50660 4678 50662 4730
rect 50662 4678 50714 4730
rect 50714 4678 50716 4730
rect 50660 4676 50716 4678
rect 50764 4730 50820 4732
rect 50764 4678 50766 4730
rect 50766 4678 50818 4730
rect 50818 4678 50820 4730
rect 50764 4676 50820 4678
rect 51996 4396 52052 4452
rect 52556 4450 52612 4452
rect 52556 4398 52558 4450
rect 52558 4398 52610 4450
rect 52610 4398 52612 4450
rect 52556 4396 52612 4398
rect 50540 4172 50596 4228
rect 50428 3500 50484 3556
rect 51884 3554 51940 3556
rect 51884 3502 51886 3554
rect 51886 3502 51938 3554
rect 51938 3502 51940 3554
rect 51884 3500 51940 3502
rect 51996 3388 52052 3444
rect 50556 3162 50612 3164
rect 50556 3110 50558 3162
rect 50558 3110 50610 3162
rect 50610 3110 50612 3162
rect 50556 3108 50612 3110
rect 50660 3162 50716 3164
rect 50660 3110 50662 3162
rect 50662 3110 50714 3162
rect 50714 3110 50716 3162
rect 50660 3108 50716 3110
rect 50764 3162 50820 3164
rect 50764 3110 50766 3162
rect 50766 3110 50818 3162
rect 50818 3110 50820 3162
rect 50764 3108 50820 3110
rect 55804 4284 55860 4340
rect 58156 45612 58212 45668
rect 58940 45666 58996 45668
rect 58940 45614 58942 45666
rect 58942 45614 58994 45666
rect 58994 45614 58996 45666
rect 58940 45612 58996 45614
rect 61292 45612 61348 45668
rect 58044 12684 58100 12740
rect 59948 14252 60004 14308
rect 65884 45724 65940 45780
rect 66556 45778 66612 45780
rect 66556 45726 66558 45778
rect 66558 45726 66610 45778
rect 66610 45726 66612 45778
rect 66556 45724 66612 45726
rect 62076 45612 62132 45668
rect 62748 45666 62804 45668
rect 62748 45614 62750 45666
rect 62750 45614 62802 45666
rect 62802 45614 62804 45666
rect 62748 45612 62804 45614
rect 69692 45612 69748 45668
rect 65916 44714 65972 44716
rect 65916 44662 65918 44714
rect 65918 44662 65970 44714
rect 65970 44662 65972 44714
rect 65916 44660 65972 44662
rect 66020 44714 66076 44716
rect 66020 44662 66022 44714
rect 66022 44662 66074 44714
rect 66074 44662 66076 44714
rect 66020 44660 66076 44662
rect 66124 44714 66180 44716
rect 66124 44662 66126 44714
rect 66126 44662 66178 44714
rect 66178 44662 66180 44714
rect 66124 44660 66180 44662
rect 65916 43146 65972 43148
rect 65916 43094 65918 43146
rect 65918 43094 65970 43146
rect 65970 43094 65972 43146
rect 65916 43092 65972 43094
rect 66020 43146 66076 43148
rect 66020 43094 66022 43146
rect 66022 43094 66074 43146
rect 66074 43094 66076 43146
rect 66020 43092 66076 43094
rect 66124 43146 66180 43148
rect 66124 43094 66126 43146
rect 66126 43094 66178 43146
rect 66178 43094 66180 43146
rect 66124 43092 66180 43094
rect 65916 41578 65972 41580
rect 65916 41526 65918 41578
rect 65918 41526 65970 41578
rect 65970 41526 65972 41578
rect 65916 41524 65972 41526
rect 66020 41578 66076 41580
rect 66020 41526 66022 41578
rect 66022 41526 66074 41578
rect 66074 41526 66076 41578
rect 66020 41524 66076 41526
rect 66124 41578 66180 41580
rect 66124 41526 66126 41578
rect 66126 41526 66178 41578
rect 66178 41526 66180 41578
rect 66124 41524 66180 41526
rect 65916 40010 65972 40012
rect 65916 39958 65918 40010
rect 65918 39958 65970 40010
rect 65970 39958 65972 40010
rect 65916 39956 65972 39958
rect 66020 40010 66076 40012
rect 66020 39958 66022 40010
rect 66022 39958 66074 40010
rect 66074 39958 66076 40010
rect 66020 39956 66076 39958
rect 66124 40010 66180 40012
rect 66124 39958 66126 40010
rect 66126 39958 66178 40010
rect 66178 39958 66180 40010
rect 66124 39956 66180 39958
rect 65916 38442 65972 38444
rect 65916 38390 65918 38442
rect 65918 38390 65970 38442
rect 65970 38390 65972 38442
rect 65916 38388 65972 38390
rect 66020 38442 66076 38444
rect 66020 38390 66022 38442
rect 66022 38390 66074 38442
rect 66074 38390 66076 38442
rect 66020 38388 66076 38390
rect 66124 38442 66180 38444
rect 66124 38390 66126 38442
rect 66126 38390 66178 38442
rect 66178 38390 66180 38442
rect 66124 38388 66180 38390
rect 65916 36874 65972 36876
rect 65916 36822 65918 36874
rect 65918 36822 65970 36874
rect 65970 36822 65972 36874
rect 65916 36820 65972 36822
rect 66020 36874 66076 36876
rect 66020 36822 66022 36874
rect 66022 36822 66074 36874
rect 66074 36822 66076 36874
rect 66020 36820 66076 36822
rect 66124 36874 66180 36876
rect 66124 36822 66126 36874
rect 66126 36822 66178 36874
rect 66178 36822 66180 36874
rect 66124 36820 66180 36822
rect 65916 35306 65972 35308
rect 65916 35254 65918 35306
rect 65918 35254 65970 35306
rect 65970 35254 65972 35306
rect 65916 35252 65972 35254
rect 66020 35306 66076 35308
rect 66020 35254 66022 35306
rect 66022 35254 66074 35306
rect 66074 35254 66076 35306
rect 66020 35252 66076 35254
rect 66124 35306 66180 35308
rect 66124 35254 66126 35306
rect 66126 35254 66178 35306
rect 66178 35254 66180 35306
rect 66124 35252 66180 35254
rect 65916 33738 65972 33740
rect 65916 33686 65918 33738
rect 65918 33686 65970 33738
rect 65970 33686 65972 33738
rect 65916 33684 65972 33686
rect 66020 33738 66076 33740
rect 66020 33686 66022 33738
rect 66022 33686 66074 33738
rect 66074 33686 66076 33738
rect 66020 33684 66076 33686
rect 66124 33738 66180 33740
rect 66124 33686 66126 33738
rect 66126 33686 66178 33738
rect 66178 33686 66180 33738
rect 66124 33684 66180 33686
rect 65916 32170 65972 32172
rect 65916 32118 65918 32170
rect 65918 32118 65970 32170
rect 65970 32118 65972 32170
rect 65916 32116 65972 32118
rect 66020 32170 66076 32172
rect 66020 32118 66022 32170
rect 66022 32118 66074 32170
rect 66074 32118 66076 32170
rect 66020 32116 66076 32118
rect 66124 32170 66180 32172
rect 66124 32118 66126 32170
rect 66126 32118 66178 32170
rect 66178 32118 66180 32170
rect 66124 32116 66180 32118
rect 65916 30602 65972 30604
rect 65916 30550 65918 30602
rect 65918 30550 65970 30602
rect 65970 30550 65972 30602
rect 65916 30548 65972 30550
rect 66020 30602 66076 30604
rect 66020 30550 66022 30602
rect 66022 30550 66074 30602
rect 66074 30550 66076 30602
rect 66020 30548 66076 30550
rect 66124 30602 66180 30604
rect 66124 30550 66126 30602
rect 66126 30550 66178 30602
rect 66178 30550 66180 30602
rect 66124 30548 66180 30550
rect 65916 29034 65972 29036
rect 65916 28982 65918 29034
rect 65918 28982 65970 29034
rect 65970 28982 65972 29034
rect 65916 28980 65972 28982
rect 66020 29034 66076 29036
rect 66020 28982 66022 29034
rect 66022 28982 66074 29034
rect 66074 28982 66076 29034
rect 66020 28980 66076 28982
rect 66124 29034 66180 29036
rect 66124 28982 66126 29034
rect 66126 28982 66178 29034
rect 66178 28982 66180 29034
rect 66124 28980 66180 28982
rect 65916 27466 65972 27468
rect 65916 27414 65918 27466
rect 65918 27414 65970 27466
rect 65970 27414 65972 27466
rect 65916 27412 65972 27414
rect 66020 27466 66076 27468
rect 66020 27414 66022 27466
rect 66022 27414 66074 27466
rect 66074 27414 66076 27466
rect 66020 27412 66076 27414
rect 66124 27466 66180 27468
rect 66124 27414 66126 27466
rect 66126 27414 66178 27466
rect 66178 27414 66180 27466
rect 66124 27412 66180 27414
rect 65916 25898 65972 25900
rect 65916 25846 65918 25898
rect 65918 25846 65970 25898
rect 65970 25846 65972 25898
rect 65916 25844 65972 25846
rect 66020 25898 66076 25900
rect 66020 25846 66022 25898
rect 66022 25846 66074 25898
rect 66074 25846 66076 25898
rect 66020 25844 66076 25846
rect 66124 25898 66180 25900
rect 66124 25846 66126 25898
rect 66126 25846 66178 25898
rect 66178 25846 66180 25898
rect 66124 25844 66180 25846
rect 65916 24330 65972 24332
rect 65916 24278 65918 24330
rect 65918 24278 65970 24330
rect 65970 24278 65972 24330
rect 65916 24276 65972 24278
rect 66020 24330 66076 24332
rect 66020 24278 66022 24330
rect 66022 24278 66074 24330
rect 66074 24278 66076 24330
rect 66020 24276 66076 24278
rect 66124 24330 66180 24332
rect 66124 24278 66126 24330
rect 66126 24278 66178 24330
rect 66178 24278 66180 24330
rect 66124 24276 66180 24278
rect 65916 22762 65972 22764
rect 65916 22710 65918 22762
rect 65918 22710 65970 22762
rect 65970 22710 65972 22762
rect 65916 22708 65972 22710
rect 66020 22762 66076 22764
rect 66020 22710 66022 22762
rect 66022 22710 66074 22762
rect 66074 22710 66076 22762
rect 66020 22708 66076 22710
rect 66124 22762 66180 22764
rect 66124 22710 66126 22762
rect 66126 22710 66178 22762
rect 66178 22710 66180 22762
rect 66124 22708 66180 22710
rect 65916 21194 65972 21196
rect 65916 21142 65918 21194
rect 65918 21142 65970 21194
rect 65970 21142 65972 21194
rect 65916 21140 65972 21142
rect 66020 21194 66076 21196
rect 66020 21142 66022 21194
rect 66022 21142 66074 21194
rect 66074 21142 66076 21194
rect 66020 21140 66076 21142
rect 66124 21194 66180 21196
rect 66124 21142 66126 21194
rect 66126 21142 66178 21194
rect 66178 21142 66180 21194
rect 66124 21140 66180 21142
rect 65916 19626 65972 19628
rect 65916 19574 65918 19626
rect 65918 19574 65970 19626
rect 65970 19574 65972 19626
rect 65916 19572 65972 19574
rect 66020 19626 66076 19628
rect 66020 19574 66022 19626
rect 66022 19574 66074 19626
rect 66074 19574 66076 19626
rect 66020 19572 66076 19574
rect 66124 19626 66180 19628
rect 66124 19574 66126 19626
rect 66126 19574 66178 19626
rect 66178 19574 66180 19626
rect 66124 19572 66180 19574
rect 68572 19292 68628 19348
rect 65916 18058 65972 18060
rect 65916 18006 65918 18058
rect 65918 18006 65970 18058
rect 65970 18006 65972 18058
rect 65916 18004 65972 18006
rect 66020 18058 66076 18060
rect 66020 18006 66022 18058
rect 66022 18006 66074 18058
rect 66074 18006 66076 18058
rect 66020 18004 66076 18006
rect 66124 18058 66180 18060
rect 66124 18006 66126 18058
rect 66126 18006 66178 18058
rect 66178 18006 66180 18058
rect 66124 18004 66180 18006
rect 65916 16490 65972 16492
rect 65916 16438 65918 16490
rect 65918 16438 65970 16490
rect 65970 16438 65972 16490
rect 65916 16436 65972 16438
rect 66020 16490 66076 16492
rect 66020 16438 66022 16490
rect 66022 16438 66074 16490
rect 66074 16438 66076 16490
rect 66020 16436 66076 16438
rect 66124 16490 66180 16492
rect 66124 16438 66126 16490
rect 66126 16438 66178 16490
rect 66178 16438 66180 16490
rect 66124 16436 66180 16438
rect 61292 14252 61348 14308
rect 63196 15932 63252 15988
rect 59948 5234 60004 5236
rect 59948 5182 59950 5234
rect 59950 5182 60002 5234
rect 60002 5182 60004 5234
rect 59948 5180 60004 5182
rect 60844 5180 60900 5236
rect 65916 14922 65972 14924
rect 65916 14870 65918 14922
rect 65918 14870 65970 14922
rect 65970 14870 65972 14922
rect 65916 14868 65972 14870
rect 66020 14922 66076 14924
rect 66020 14870 66022 14922
rect 66022 14870 66074 14922
rect 66074 14870 66076 14922
rect 66020 14868 66076 14870
rect 66124 14922 66180 14924
rect 66124 14870 66126 14922
rect 66126 14870 66178 14922
rect 66178 14870 66180 14922
rect 66124 14868 66180 14870
rect 65916 13354 65972 13356
rect 65916 13302 65918 13354
rect 65918 13302 65970 13354
rect 65970 13302 65972 13354
rect 65916 13300 65972 13302
rect 66020 13354 66076 13356
rect 66020 13302 66022 13354
rect 66022 13302 66074 13354
rect 66074 13302 66076 13354
rect 66020 13300 66076 13302
rect 66124 13354 66180 13356
rect 66124 13302 66126 13354
rect 66126 13302 66178 13354
rect 66178 13302 66180 13354
rect 66124 13300 66180 13302
rect 65916 11786 65972 11788
rect 65916 11734 65918 11786
rect 65918 11734 65970 11786
rect 65970 11734 65972 11786
rect 65916 11732 65972 11734
rect 66020 11786 66076 11788
rect 66020 11734 66022 11786
rect 66022 11734 66074 11786
rect 66074 11734 66076 11786
rect 66020 11732 66076 11734
rect 66124 11786 66180 11788
rect 66124 11734 66126 11786
rect 66126 11734 66178 11786
rect 66178 11734 66180 11786
rect 66124 11732 66180 11734
rect 65436 11228 65492 11284
rect 65916 10218 65972 10220
rect 65916 10166 65918 10218
rect 65918 10166 65970 10218
rect 65970 10166 65972 10218
rect 65916 10164 65972 10166
rect 66020 10218 66076 10220
rect 66020 10166 66022 10218
rect 66022 10166 66074 10218
rect 66074 10166 66076 10218
rect 66020 10164 66076 10166
rect 66124 10218 66180 10220
rect 66124 10166 66126 10218
rect 66126 10166 66178 10218
rect 66178 10166 66180 10218
rect 66124 10164 66180 10166
rect 65916 8650 65972 8652
rect 65916 8598 65918 8650
rect 65918 8598 65970 8650
rect 65970 8598 65972 8650
rect 65916 8596 65972 8598
rect 66020 8650 66076 8652
rect 66020 8598 66022 8650
rect 66022 8598 66074 8650
rect 66074 8598 66076 8650
rect 66020 8596 66076 8598
rect 66124 8650 66180 8652
rect 66124 8598 66126 8650
rect 66126 8598 66178 8650
rect 66178 8598 66180 8650
rect 66124 8596 66180 8598
rect 65916 7082 65972 7084
rect 65916 7030 65918 7082
rect 65918 7030 65970 7082
rect 65970 7030 65972 7082
rect 65916 7028 65972 7030
rect 66020 7082 66076 7084
rect 66020 7030 66022 7082
rect 66022 7030 66074 7082
rect 66074 7030 66076 7082
rect 66020 7028 66076 7030
rect 66124 7082 66180 7084
rect 66124 7030 66126 7082
rect 66126 7030 66178 7082
rect 66178 7030 66180 7082
rect 66124 7028 66180 7030
rect 65916 5514 65972 5516
rect 65916 5462 65918 5514
rect 65918 5462 65970 5514
rect 65970 5462 65972 5514
rect 65916 5460 65972 5462
rect 66020 5514 66076 5516
rect 66020 5462 66022 5514
rect 66022 5462 66074 5514
rect 66074 5462 66076 5514
rect 66020 5460 66076 5462
rect 66124 5514 66180 5516
rect 66124 5462 66126 5514
rect 66126 5462 66178 5514
rect 66178 5462 66180 5514
rect 66124 5460 66180 5462
rect 69916 45612 69972 45668
rect 70364 45666 70420 45668
rect 70364 45614 70366 45666
rect 70366 45614 70418 45666
rect 70418 45614 70420 45666
rect 70364 45612 70420 45614
rect 73276 45612 73332 45668
rect 73500 45612 73556 45668
rect 74172 45666 74228 45668
rect 74172 45614 74174 45666
rect 74174 45614 74226 45666
rect 74226 45614 74228 45666
rect 74172 45612 74228 45614
rect 96636 46282 96692 46284
rect 96636 46230 96638 46282
rect 96638 46230 96690 46282
rect 96690 46230 96692 46282
rect 96636 46228 96692 46230
rect 96740 46282 96796 46284
rect 96740 46230 96742 46282
rect 96742 46230 96794 46282
rect 96794 46230 96796 46282
rect 96740 46228 96796 46230
rect 96844 46282 96900 46284
rect 96844 46230 96846 46282
rect 96846 46230 96898 46282
rect 96898 46230 96900 46282
rect 96844 46228 96900 46230
rect 100156 45836 100212 45892
rect 100828 45890 100884 45892
rect 100828 45838 100830 45890
rect 100830 45838 100882 45890
rect 100882 45838 100884 45890
rect 100828 45836 100884 45838
rect 103964 45836 104020 45892
rect 104636 45890 104692 45892
rect 104636 45838 104638 45890
rect 104638 45838 104690 45890
rect 104690 45838 104692 45890
rect 104636 45836 104692 45838
rect 127356 46282 127412 46284
rect 127356 46230 127358 46282
rect 127358 46230 127410 46282
rect 127410 46230 127412 46282
rect 127356 46228 127412 46230
rect 127460 46282 127516 46284
rect 127460 46230 127462 46282
rect 127462 46230 127514 46282
rect 127514 46230 127516 46282
rect 127460 46228 127516 46230
rect 127564 46282 127620 46284
rect 127564 46230 127566 46282
rect 127566 46230 127618 46282
rect 127618 46230 127620 46282
rect 127564 46228 127620 46230
rect 148092 46060 148148 46116
rect 150444 46114 150500 46116
rect 150444 46062 150446 46114
rect 150446 46062 150498 46114
rect 150498 46062 150500 46114
rect 150444 46060 150500 46062
rect 150332 45948 150388 46004
rect 130172 45724 130228 45780
rect 76412 45612 76468 45668
rect 81276 45498 81332 45500
rect 81276 45446 81278 45498
rect 81278 45446 81330 45498
rect 81330 45446 81332 45498
rect 81276 45444 81332 45446
rect 81380 45498 81436 45500
rect 81380 45446 81382 45498
rect 81382 45446 81434 45498
rect 81434 45446 81436 45498
rect 81380 45444 81436 45446
rect 81484 45498 81540 45500
rect 81484 45446 81486 45498
rect 81486 45446 81538 45498
rect 81538 45446 81540 45498
rect 81484 45444 81540 45446
rect 81276 43930 81332 43932
rect 81276 43878 81278 43930
rect 81278 43878 81330 43930
rect 81330 43878 81332 43930
rect 81276 43876 81332 43878
rect 81380 43930 81436 43932
rect 81380 43878 81382 43930
rect 81382 43878 81434 43930
rect 81434 43878 81436 43930
rect 81380 43876 81436 43878
rect 81484 43930 81540 43932
rect 81484 43878 81486 43930
rect 81486 43878 81538 43930
rect 81538 43878 81540 43930
rect 81484 43876 81540 43878
rect 80108 43596 80164 43652
rect 81276 42362 81332 42364
rect 81276 42310 81278 42362
rect 81278 42310 81330 42362
rect 81330 42310 81332 42362
rect 81276 42308 81332 42310
rect 81380 42362 81436 42364
rect 81380 42310 81382 42362
rect 81382 42310 81434 42362
rect 81434 42310 81436 42362
rect 81380 42308 81436 42310
rect 81484 42362 81540 42364
rect 81484 42310 81486 42362
rect 81486 42310 81538 42362
rect 81538 42310 81540 42362
rect 81484 42308 81540 42310
rect 81276 40794 81332 40796
rect 81276 40742 81278 40794
rect 81278 40742 81330 40794
rect 81330 40742 81332 40794
rect 81276 40740 81332 40742
rect 81380 40794 81436 40796
rect 81380 40742 81382 40794
rect 81382 40742 81434 40794
rect 81434 40742 81436 40794
rect 81380 40740 81436 40742
rect 81484 40794 81540 40796
rect 81484 40742 81486 40794
rect 81486 40742 81538 40794
rect 81538 40742 81540 40794
rect 81484 40740 81540 40742
rect 81276 39226 81332 39228
rect 81276 39174 81278 39226
rect 81278 39174 81330 39226
rect 81330 39174 81332 39226
rect 81276 39172 81332 39174
rect 81380 39226 81436 39228
rect 81380 39174 81382 39226
rect 81382 39174 81434 39226
rect 81434 39174 81436 39226
rect 81380 39172 81436 39174
rect 81484 39226 81540 39228
rect 81484 39174 81486 39226
rect 81486 39174 81538 39226
rect 81538 39174 81540 39226
rect 81484 39172 81540 39174
rect 81276 37658 81332 37660
rect 81276 37606 81278 37658
rect 81278 37606 81330 37658
rect 81330 37606 81332 37658
rect 81276 37604 81332 37606
rect 81380 37658 81436 37660
rect 81380 37606 81382 37658
rect 81382 37606 81434 37658
rect 81434 37606 81436 37658
rect 81380 37604 81436 37606
rect 81484 37658 81540 37660
rect 81484 37606 81486 37658
rect 81486 37606 81538 37658
rect 81538 37606 81540 37658
rect 81484 37604 81540 37606
rect 81276 36090 81332 36092
rect 81276 36038 81278 36090
rect 81278 36038 81330 36090
rect 81330 36038 81332 36090
rect 81276 36036 81332 36038
rect 81380 36090 81436 36092
rect 81380 36038 81382 36090
rect 81382 36038 81434 36090
rect 81434 36038 81436 36090
rect 81380 36036 81436 36038
rect 81484 36090 81540 36092
rect 81484 36038 81486 36090
rect 81486 36038 81538 36090
rect 81538 36038 81540 36090
rect 81484 36036 81540 36038
rect 96636 44714 96692 44716
rect 96636 44662 96638 44714
rect 96638 44662 96690 44714
rect 96690 44662 96692 44714
rect 96636 44660 96692 44662
rect 96740 44714 96796 44716
rect 96740 44662 96742 44714
rect 96742 44662 96794 44714
rect 96794 44662 96796 44714
rect 96740 44660 96796 44662
rect 96844 44714 96900 44716
rect 96844 44662 96846 44714
rect 96846 44662 96898 44714
rect 96898 44662 96900 44714
rect 96844 44660 96900 44662
rect 96636 43146 96692 43148
rect 96636 43094 96638 43146
rect 96638 43094 96690 43146
rect 96690 43094 96692 43146
rect 96636 43092 96692 43094
rect 96740 43146 96796 43148
rect 96740 43094 96742 43146
rect 96742 43094 96794 43146
rect 96794 43094 96796 43146
rect 96740 43092 96796 43094
rect 96844 43146 96900 43148
rect 96844 43094 96846 43146
rect 96846 43094 96898 43146
rect 96898 43094 96900 43146
rect 96844 43092 96900 43094
rect 96636 41578 96692 41580
rect 96636 41526 96638 41578
rect 96638 41526 96690 41578
rect 96690 41526 96692 41578
rect 96636 41524 96692 41526
rect 96740 41578 96796 41580
rect 96740 41526 96742 41578
rect 96742 41526 96794 41578
rect 96794 41526 96796 41578
rect 96740 41524 96796 41526
rect 96844 41578 96900 41580
rect 96844 41526 96846 41578
rect 96846 41526 96898 41578
rect 96898 41526 96900 41578
rect 96844 41524 96900 41526
rect 92204 41132 92260 41188
rect 96636 40010 96692 40012
rect 96636 39958 96638 40010
rect 96638 39958 96690 40010
rect 96690 39958 96692 40010
rect 96636 39956 96692 39958
rect 96740 40010 96796 40012
rect 96740 39958 96742 40010
rect 96742 39958 96794 40010
rect 96794 39958 96796 40010
rect 96740 39956 96796 39958
rect 96844 40010 96900 40012
rect 96844 39958 96846 40010
rect 96846 39958 96898 40010
rect 96898 39958 96900 40010
rect 96844 39956 96900 39958
rect 88172 39452 88228 39508
rect 96636 38442 96692 38444
rect 96636 38390 96638 38442
rect 96638 38390 96690 38442
rect 96690 38390 96692 38442
rect 96636 38388 96692 38390
rect 96740 38442 96796 38444
rect 96740 38390 96742 38442
rect 96742 38390 96794 38442
rect 96794 38390 96796 38442
rect 96740 38388 96796 38390
rect 96844 38442 96900 38444
rect 96844 38390 96846 38442
rect 96846 38390 96898 38442
rect 96898 38390 96900 38442
rect 96844 38388 96900 38390
rect 96636 36874 96692 36876
rect 96636 36822 96638 36874
rect 96638 36822 96690 36874
rect 96690 36822 96692 36874
rect 96636 36820 96692 36822
rect 96740 36874 96796 36876
rect 96740 36822 96742 36874
rect 96742 36822 96794 36874
rect 96794 36822 96796 36874
rect 96740 36820 96796 36822
rect 96844 36874 96900 36876
rect 96844 36822 96846 36874
rect 96846 36822 96898 36874
rect 96898 36822 96900 36874
rect 96844 36820 96900 36822
rect 96636 35306 96692 35308
rect 96636 35254 96638 35306
rect 96638 35254 96690 35306
rect 96690 35254 96692 35306
rect 96636 35252 96692 35254
rect 96740 35306 96796 35308
rect 96740 35254 96742 35306
rect 96742 35254 96794 35306
rect 96794 35254 96796 35306
rect 96740 35252 96796 35254
rect 96844 35306 96900 35308
rect 96844 35254 96846 35306
rect 96846 35254 96898 35306
rect 96898 35254 96900 35306
rect 96844 35252 96900 35254
rect 84140 34636 84196 34692
rect 81276 34522 81332 34524
rect 81276 34470 81278 34522
rect 81278 34470 81330 34522
rect 81330 34470 81332 34522
rect 81276 34468 81332 34470
rect 81380 34522 81436 34524
rect 81380 34470 81382 34522
rect 81382 34470 81434 34522
rect 81434 34470 81436 34522
rect 81380 34468 81436 34470
rect 81484 34522 81540 34524
rect 81484 34470 81486 34522
rect 81486 34470 81538 34522
rect 81538 34470 81540 34522
rect 81484 34468 81540 34470
rect 96636 33738 96692 33740
rect 96636 33686 96638 33738
rect 96638 33686 96690 33738
rect 96690 33686 96692 33738
rect 96636 33684 96692 33686
rect 96740 33738 96796 33740
rect 96740 33686 96742 33738
rect 96742 33686 96794 33738
rect 96794 33686 96796 33738
rect 96740 33684 96796 33686
rect 96844 33738 96900 33740
rect 96844 33686 96846 33738
rect 96846 33686 96898 33738
rect 96898 33686 96900 33738
rect 96844 33684 96900 33686
rect 81276 32954 81332 32956
rect 81276 32902 81278 32954
rect 81278 32902 81330 32954
rect 81330 32902 81332 32954
rect 81276 32900 81332 32902
rect 81380 32954 81436 32956
rect 81380 32902 81382 32954
rect 81382 32902 81434 32954
rect 81434 32902 81436 32954
rect 81380 32900 81436 32902
rect 81484 32954 81540 32956
rect 81484 32902 81486 32954
rect 81486 32902 81538 32954
rect 81538 32902 81540 32954
rect 81484 32900 81540 32902
rect 96636 32170 96692 32172
rect 96636 32118 96638 32170
rect 96638 32118 96690 32170
rect 96690 32118 96692 32170
rect 96636 32116 96692 32118
rect 96740 32170 96796 32172
rect 96740 32118 96742 32170
rect 96742 32118 96794 32170
rect 96794 32118 96796 32170
rect 96740 32116 96796 32118
rect 96844 32170 96900 32172
rect 96844 32118 96846 32170
rect 96846 32118 96898 32170
rect 96898 32118 96900 32170
rect 96844 32116 96900 32118
rect 76412 19292 76468 19348
rect 73276 17612 73332 17668
rect 69692 15932 69748 15988
rect 81276 31386 81332 31388
rect 81276 31334 81278 31386
rect 81278 31334 81330 31386
rect 81330 31334 81332 31386
rect 81276 31332 81332 31334
rect 81380 31386 81436 31388
rect 81380 31334 81382 31386
rect 81382 31334 81434 31386
rect 81434 31334 81436 31386
rect 81380 31332 81436 31334
rect 81484 31386 81540 31388
rect 81484 31334 81486 31386
rect 81486 31334 81538 31386
rect 81538 31334 81540 31386
rect 81484 31332 81540 31334
rect 96636 30602 96692 30604
rect 96636 30550 96638 30602
rect 96638 30550 96690 30602
rect 96690 30550 96692 30602
rect 96636 30548 96692 30550
rect 96740 30602 96796 30604
rect 96740 30550 96742 30602
rect 96742 30550 96794 30602
rect 96794 30550 96796 30602
rect 96740 30548 96796 30550
rect 96844 30602 96900 30604
rect 96844 30550 96846 30602
rect 96846 30550 96898 30602
rect 96898 30550 96900 30602
rect 96844 30548 96900 30550
rect 96236 30210 96292 30212
rect 96236 30158 96238 30210
rect 96238 30158 96290 30210
rect 96290 30158 96292 30210
rect 96236 30156 96292 30158
rect 96684 30210 96740 30212
rect 96684 30158 96686 30210
rect 96686 30158 96738 30210
rect 96738 30158 96740 30210
rect 96684 30156 96740 30158
rect 93772 30044 93828 30100
rect 81276 29818 81332 29820
rect 81276 29766 81278 29818
rect 81278 29766 81330 29818
rect 81330 29766 81332 29818
rect 81276 29764 81332 29766
rect 81380 29818 81436 29820
rect 81380 29766 81382 29818
rect 81382 29766 81434 29818
rect 81434 29766 81436 29818
rect 81380 29764 81436 29766
rect 81484 29818 81540 29820
rect 81484 29766 81486 29818
rect 81486 29766 81538 29818
rect 81538 29766 81540 29818
rect 81484 29764 81540 29766
rect 81276 28250 81332 28252
rect 81276 28198 81278 28250
rect 81278 28198 81330 28250
rect 81330 28198 81332 28250
rect 81276 28196 81332 28198
rect 81380 28250 81436 28252
rect 81380 28198 81382 28250
rect 81382 28198 81434 28250
rect 81434 28198 81436 28250
rect 81380 28196 81436 28198
rect 81484 28250 81540 28252
rect 81484 28198 81486 28250
rect 81486 28198 81538 28250
rect 81538 28198 81540 28250
rect 81484 28196 81540 28198
rect 81276 26682 81332 26684
rect 81276 26630 81278 26682
rect 81278 26630 81330 26682
rect 81330 26630 81332 26682
rect 81276 26628 81332 26630
rect 81380 26682 81436 26684
rect 81380 26630 81382 26682
rect 81382 26630 81434 26682
rect 81434 26630 81436 26682
rect 81380 26628 81436 26630
rect 81484 26682 81540 26684
rect 81484 26630 81486 26682
rect 81486 26630 81538 26682
rect 81538 26630 81540 26682
rect 81484 26628 81540 26630
rect 81276 25114 81332 25116
rect 81276 25062 81278 25114
rect 81278 25062 81330 25114
rect 81330 25062 81332 25114
rect 81276 25060 81332 25062
rect 81380 25114 81436 25116
rect 81380 25062 81382 25114
rect 81382 25062 81434 25114
rect 81434 25062 81436 25114
rect 81380 25060 81436 25062
rect 81484 25114 81540 25116
rect 81484 25062 81486 25114
rect 81486 25062 81538 25114
rect 81538 25062 81540 25114
rect 81484 25060 81540 25062
rect 81276 23546 81332 23548
rect 81276 23494 81278 23546
rect 81278 23494 81330 23546
rect 81330 23494 81332 23546
rect 81276 23492 81332 23494
rect 81380 23546 81436 23548
rect 81380 23494 81382 23546
rect 81382 23494 81434 23546
rect 81434 23494 81436 23546
rect 81380 23492 81436 23494
rect 81484 23546 81540 23548
rect 81484 23494 81486 23546
rect 81486 23494 81538 23546
rect 81538 23494 81540 23546
rect 81484 23492 81540 23494
rect 81276 21978 81332 21980
rect 81276 21926 81278 21978
rect 81278 21926 81330 21978
rect 81330 21926 81332 21978
rect 81276 21924 81332 21926
rect 81380 21978 81436 21980
rect 81380 21926 81382 21978
rect 81382 21926 81434 21978
rect 81434 21926 81436 21978
rect 81380 21924 81436 21926
rect 81484 21978 81540 21980
rect 81484 21926 81486 21978
rect 81486 21926 81538 21978
rect 81538 21926 81540 21978
rect 81484 21924 81540 21926
rect 81276 20410 81332 20412
rect 81276 20358 81278 20410
rect 81278 20358 81330 20410
rect 81330 20358 81332 20410
rect 81276 20356 81332 20358
rect 81380 20410 81436 20412
rect 81380 20358 81382 20410
rect 81382 20358 81434 20410
rect 81434 20358 81436 20410
rect 81380 20356 81436 20358
rect 81484 20410 81540 20412
rect 81484 20358 81486 20410
rect 81486 20358 81538 20410
rect 81538 20358 81540 20410
rect 81484 20356 81540 20358
rect 81276 18842 81332 18844
rect 81276 18790 81278 18842
rect 81278 18790 81330 18842
rect 81330 18790 81332 18842
rect 81276 18788 81332 18790
rect 81380 18842 81436 18844
rect 81380 18790 81382 18842
rect 81382 18790 81434 18842
rect 81434 18790 81436 18842
rect 81380 18788 81436 18790
rect 81484 18842 81540 18844
rect 81484 18790 81486 18842
rect 81486 18790 81538 18842
rect 81538 18790 81540 18842
rect 81484 18788 81540 18790
rect 81276 17274 81332 17276
rect 81276 17222 81278 17274
rect 81278 17222 81330 17274
rect 81330 17222 81332 17274
rect 81276 17220 81332 17222
rect 81380 17274 81436 17276
rect 81380 17222 81382 17274
rect 81382 17222 81434 17274
rect 81434 17222 81436 17274
rect 81380 17220 81436 17222
rect 81484 17274 81540 17276
rect 81484 17222 81486 17274
rect 81486 17222 81538 17274
rect 81538 17222 81540 17274
rect 81484 17220 81540 17222
rect 81276 15706 81332 15708
rect 81276 15654 81278 15706
rect 81278 15654 81330 15706
rect 81330 15654 81332 15706
rect 81276 15652 81332 15654
rect 81380 15706 81436 15708
rect 81380 15654 81382 15706
rect 81382 15654 81434 15706
rect 81434 15654 81436 15706
rect 81380 15652 81436 15654
rect 81484 15706 81540 15708
rect 81484 15654 81486 15706
rect 81486 15654 81538 15706
rect 81538 15654 81540 15706
rect 81484 15652 81540 15654
rect 81276 14138 81332 14140
rect 81276 14086 81278 14138
rect 81278 14086 81330 14138
rect 81330 14086 81332 14138
rect 81276 14084 81332 14086
rect 81380 14138 81436 14140
rect 81380 14086 81382 14138
rect 81382 14086 81434 14138
rect 81434 14086 81436 14138
rect 81380 14084 81436 14086
rect 81484 14138 81540 14140
rect 81484 14086 81486 14138
rect 81486 14086 81538 14138
rect 81538 14086 81540 14138
rect 81484 14084 81540 14086
rect 81276 12570 81332 12572
rect 81276 12518 81278 12570
rect 81278 12518 81330 12570
rect 81330 12518 81332 12570
rect 81276 12516 81332 12518
rect 81380 12570 81436 12572
rect 81380 12518 81382 12570
rect 81382 12518 81434 12570
rect 81434 12518 81436 12570
rect 81380 12516 81436 12518
rect 81484 12570 81540 12572
rect 81484 12518 81486 12570
rect 81486 12518 81538 12570
rect 81538 12518 81540 12570
rect 81484 12516 81540 12518
rect 77868 11228 77924 11284
rect 81276 11002 81332 11004
rect 81276 10950 81278 11002
rect 81278 10950 81330 11002
rect 81330 10950 81332 11002
rect 81276 10948 81332 10950
rect 81380 11002 81436 11004
rect 81380 10950 81382 11002
rect 81382 10950 81434 11002
rect 81434 10950 81436 11002
rect 81380 10948 81436 10950
rect 81484 11002 81540 11004
rect 81484 10950 81486 11002
rect 81486 10950 81538 11002
rect 81538 10950 81540 11002
rect 81484 10948 81540 10950
rect 81276 9434 81332 9436
rect 81276 9382 81278 9434
rect 81278 9382 81330 9434
rect 81330 9382 81332 9434
rect 81276 9380 81332 9382
rect 81380 9434 81436 9436
rect 81380 9382 81382 9434
rect 81382 9382 81434 9434
rect 81434 9382 81436 9434
rect 81380 9380 81436 9382
rect 81484 9434 81540 9436
rect 81484 9382 81486 9434
rect 81486 9382 81538 9434
rect 81538 9382 81540 9434
rect 81484 9380 81540 9382
rect 88060 8428 88116 8484
rect 81276 7866 81332 7868
rect 81276 7814 81278 7866
rect 81278 7814 81330 7866
rect 81330 7814 81332 7866
rect 81276 7812 81332 7814
rect 81380 7866 81436 7868
rect 81380 7814 81382 7866
rect 81382 7814 81434 7866
rect 81434 7814 81436 7866
rect 81380 7812 81436 7814
rect 81484 7866 81540 7868
rect 81484 7814 81486 7866
rect 81486 7814 81538 7866
rect 81538 7814 81540 7866
rect 81484 7812 81540 7814
rect 73052 6412 73108 6468
rect 57596 4338 57652 4340
rect 57596 4286 57598 4338
rect 57598 4286 57650 4338
rect 57650 4286 57652 4338
rect 57596 4284 57652 4286
rect 57036 4172 57092 4228
rect 57372 4060 57428 4116
rect 56028 3666 56084 3668
rect 56028 3614 56030 3666
rect 56030 3614 56082 3666
rect 56082 3614 56084 3666
rect 56028 3612 56084 3614
rect 53116 3500 53172 3556
rect 55020 3554 55076 3556
rect 55020 3502 55022 3554
rect 55022 3502 55074 3554
rect 55074 3502 55076 3554
rect 55020 3500 55076 3502
rect 52892 3388 52948 3444
rect 54684 3388 54740 3444
rect 58604 4114 58660 4116
rect 58604 4062 58606 4114
rect 58606 4062 58658 4114
rect 58658 4062 58660 4114
rect 58604 4060 58660 4062
rect 58492 3500 58548 3556
rect 59500 3554 59556 3556
rect 59500 3502 59502 3554
rect 59502 3502 59554 3554
rect 59554 3502 59556 3554
rect 59500 3500 59556 3502
rect 61180 3500 61236 3556
rect 62748 3612 62804 3668
rect 62972 3554 63028 3556
rect 62972 3502 62974 3554
rect 62974 3502 63026 3554
rect 63026 3502 63028 3554
rect 62972 3500 63028 3502
rect 66556 4284 66612 4340
rect 68348 4338 68404 4340
rect 68348 4286 68350 4338
rect 68350 4286 68402 4338
rect 68402 4286 68404 4338
rect 68348 4284 68404 4286
rect 68124 4060 68180 4116
rect 65916 3946 65972 3948
rect 65916 3894 65918 3946
rect 65918 3894 65970 3946
rect 65970 3894 65972 3946
rect 65916 3892 65972 3894
rect 66020 3946 66076 3948
rect 66020 3894 66022 3946
rect 66022 3894 66074 3946
rect 66074 3894 66076 3946
rect 66020 3892 66076 3894
rect 66124 3946 66180 3948
rect 66124 3894 66126 3946
rect 66126 3894 66178 3946
rect 66178 3894 66180 3946
rect 66124 3892 66180 3894
rect 63980 3666 64036 3668
rect 63980 3614 63982 3666
rect 63982 3614 64034 3666
rect 64034 3614 64036 3666
rect 63980 3612 64036 3614
rect 67452 3666 67508 3668
rect 67452 3614 67454 3666
rect 67454 3614 67506 3666
rect 67506 3614 67508 3666
rect 67452 3612 67508 3614
rect 63868 3500 63924 3556
rect 66444 3554 66500 3556
rect 66444 3502 66446 3554
rect 66446 3502 66498 3554
rect 66498 3502 66500 3554
rect 66444 3500 66500 3502
rect 65436 3388 65492 3444
rect 81276 6298 81332 6300
rect 81276 6246 81278 6298
rect 81278 6246 81330 6298
rect 81330 6246 81332 6298
rect 81276 6244 81332 6246
rect 81380 6298 81436 6300
rect 81380 6246 81382 6298
rect 81382 6246 81434 6298
rect 81434 6246 81436 6298
rect 81380 6244 81436 6246
rect 81484 6298 81540 6300
rect 81484 6246 81486 6298
rect 81486 6246 81538 6298
rect 81538 6246 81540 6298
rect 81484 6244 81540 6246
rect 84252 5628 84308 5684
rect 81276 4730 81332 4732
rect 81276 4678 81278 4730
rect 81278 4678 81330 4730
rect 81330 4678 81332 4730
rect 81276 4676 81332 4678
rect 81380 4730 81436 4732
rect 81380 4678 81382 4730
rect 81382 4678 81434 4730
rect 81434 4678 81436 4730
rect 81380 4676 81436 4678
rect 81484 4730 81540 4732
rect 81484 4678 81486 4730
rect 81486 4678 81538 4730
rect 81538 4678 81540 4730
rect 81484 4676 81540 4678
rect 73052 4396 73108 4452
rect 77196 4396 77252 4452
rect 69356 4114 69412 4116
rect 69356 4062 69358 4114
rect 69358 4062 69410 4114
rect 69410 4062 69412 4114
rect 69356 4060 69412 4062
rect 73500 3612 73556 3668
rect 69244 3500 69300 3556
rect 70924 3554 70980 3556
rect 70924 3502 70926 3554
rect 70926 3502 70978 3554
rect 70978 3502 70980 3554
rect 70924 3500 70980 3502
rect 70812 3388 70868 3444
rect 71932 3388 71988 3444
rect 74284 3666 74340 3668
rect 74284 3614 74286 3666
rect 74286 3614 74338 3666
rect 74338 3614 74340 3666
rect 74284 3612 74340 3614
rect 76524 3612 76580 3668
rect 78876 4338 78932 4340
rect 78876 4286 78878 4338
rect 78878 4286 78930 4338
rect 78930 4286 78932 4338
rect 78876 4284 78932 4286
rect 79548 4338 79604 4340
rect 79548 4286 79550 4338
rect 79550 4286 79602 4338
rect 79602 4286 79604 4338
rect 79548 4284 79604 4286
rect 80556 4284 80612 4340
rect 77196 3666 77252 3668
rect 77196 3614 77198 3666
rect 77198 3614 77250 3666
rect 77250 3614 77252 3666
rect 77196 3612 77252 3614
rect 81340 4338 81396 4340
rect 81340 4286 81342 4338
rect 81342 4286 81394 4338
rect 81394 4286 81396 4338
rect 81340 4284 81396 4286
rect 92764 5740 92820 5796
rect 89068 5292 89124 5348
rect 95452 30098 95508 30100
rect 95452 30046 95454 30098
rect 95454 30046 95506 30098
rect 95506 30046 95508 30098
rect 95452 30044 95508 30046
rect 97132 30098 97188 30100
rect 97132 30046 97134 30098
rect 97134 30046 97186 30098
rect 97186 30046 97188 30098
rect 97132 30044 97188 30046
rect 101276 30156 101332 30212
rect 101612 30044 101668 30100
rect 97916 29260 97972 29316
rect 96636 29034 96692 29036
rect 96636 28982 96638 29034
rect 96638 28982 96690 29034
rect 96690 28982 96692 29034
rect 96636 28980 96692 28982
rect 96740 29034 96796 29036
rect 96740 28982 96742 29034
rect 96742 28982 96794 29034
rect 96794 28982 96796 29034
rect 96740 28980 96796 28982
rect 96844 29034 96900 29036
rect 96844 28982 96846 29034
rect 96846 28982 96898 29034
rect 96898 28982 96900 29034
rect 96844 28980 96900 28982
rect 96636 27466 96692 27468
rect 96636 27414 96638 27466
rect 96638 27414 96690 27466
rect 96690 27414 96692 27466
rect 96636 27412 96692 27414
rect 96740 27466 96796 27468
rect 96740 27414 96742 27466
rect 96742 27414 96794 27466
rect 96794 27414 96796 27466
rect 96740 27412 96796 27414
rect 96844 27466 96900 27468
rect 96844 27414 96846 27466
rect 96846 27414 96898 27466
rect 96898 27414 96900 27466
rect 96844 27412 96900 27414
rect 96636 25898 96692 25900
rect 96636 25846 96638 25898
rect 96638 25846 96690 25898
rect 96690 25846 96692 25898
rect 96636 25844 96692 25846
rect 96740 25898 96796 25900
rect 96740 25846 96742 25898
rect 96742 25846 96794 25898
rect 96794 25846 96796 25898
rect 96740 25844 96796 25846
rect 96844 25898 96900 25900
rect 96844 25846 96846 25898
rect 96846 25846 96898 25898
rect 96898 25846 96900 25898
rect 96844 25844 96900 25846
rect 96636 24330 96692 24332
rect 96636 24278 96638 24330
rect 96638 24278 96690 24330
rect 96690 24278 96692 24330
rect 96636 24276 96692 24278
rect 96740 24330 96796 24332
rect 96740 24278 96742 24330
rect 96742 24278 96794 24330
rect 96794 24278 96796 24330
rect 96740 24276 96796 24278
rect 96844 24330 96900 24332
rect 96844 24278 96846 24330
rect 96846 24278 96898 24330
rect 96898 24278 96900 24330
rect 96844 24276 96900 24278
rect 96636 22762 96692 22764
rect 96636 22710 96638 22762
rect 96638 22710 96690 22762
rect 96690 22710 96692 22762
rect 96636 22708 96692 22710
rect 96740 22762 96796 22764
rect 96740 22710 96742 22762
rect 96742 22710 96794 22762
rect 96794 22710 96796 22762
rect 96740 22708 96796 22710
rect 96844 22762 96900 22764
rect 96844 22710 96846 22762
rect 96846 22710 96898 22762
rect 96898 22710 96900 22762
rect 96844 22708 96900 22710
rect 96636 21194 96692 21196
rect 96636 21142 96638 21194
rect 96638 21142 96690 21194
rect 96690 21142 96692 21194
rect 96636 21140 96692 21142
rect 96740 21194 96796 21196
rect 96740 21142 96742 21194
rect 96742 21142 96794 21194
rect 96794 21142 96796 21194
rect 96740 21140 96796 21142
rect 96844 21194 96900 21196
rect 96844 21142 96846 21194
rect 96846 21142 96898 21194
rect 96898 21142 96900 21194
rect 96844 21140 96900 21142
rect 96636 19626 96692 19628
rect 96636 19574 96638 19626
rect 96638 19574 96690 19626
rect 96690 19574 96692 19626
rect 96636 19572 96692 19574
rect 96740 19626 96796 19628
rect 96740 19574 96742 19626
rect 96742 19574 96794 19626
rect 96794 19574 96796 19626
rect 96740 19572 96796 19574
rect 96844 19626 96900 19628
rect 96844 19574 96846 19626
rect 96846 19574 96898 19626
rect 96898 19574 96900 19626
rect 96844 19572 96900 19574
rect 96636 18058 96692 18060
rect 96636 18006 96638 18058
rect 96638 18006 96690 18058
rect 96690 18006 96692 18058
rect 96636 18004 96692 18006
rect 96740 18058 96796 18060
rect 96740 18006 96742 18058
rect 96742 18006 96794 18058
rect 96794 18006 96796 18058
rect 96740 18004 96796 18006
rect 96844 18058 96900 18060
rect 96844 18006 96846 18058
rect 96846 18006 96898 18058
rect 96898 18006 96900 18058
rect 96844 18004 96900 18006
rect 96636 16490 96692 16492
rect 96636 16438 96638 16490
rect 96638 16438 96690 16490
rect 96690 16438 96692 16490
rect 96636 16436 96692 16438
rect 96740 16490 96796 16492
rect 96740 16438 96742 16490
rect 96742 16438 96794 16490
rect 96794 16438 96796 16490
rect 96740 16436 96796 16438
rect 96844 16490 96900 16492
rect 96844 16438 96846 16490
rect 96846 16438 96898 16490
rect 96898 16438 96900 16490
rect 96844 16436 96900 16438
rect 96636 14922 96692 14924
rect 96636 14870 96638 14922
rect 96638 14870 96690 14922
rect 96690 14870 96692 14922
rect 96636 14868 96692 14870
rect 96740 14922 96796 14924
rect 96740 14870 96742 14922
rect 96742 14870 96794 14922
rect 96794 14870 96796 14922
rect 96740 14868 96796 14870
rect 96844 14922 96900 14924
rect 96844 14870 96846 14922
rect 96846 14870 96898 14922
rect 96898 14870 96900 14922
rect 96844 14868 96900 14870
rect 96636 13354 96692 13356
rect 96636 13302 96638 13354
rect 96638 13302 96690 13354
rect 96690 13302 96692 13354
rect 96636 13300 96692 13302
rect 96740 13354 96796 13356
rect 96740 13302 96742 13354
rect 96742 13302 96794 13354
rect 96794 13302 96796 13354
rect 96740 13300 96796 13302
rect 96844 13354 96900 13356
rect 96844 13302 96846 13354
rect 96846 13302 96898 13354
rect 96898 13302 96900 13354
rect 96844 13300 96900 13302
rect 96636 11786 96692 11788
rect 96636 11734 96638 11786
rect 96638 11734 96690 11786
rect 96690 11734 96692 11786
rect 96636 11732 96692 11734
rect 96740 11786 96796 11788
rect 96740 11734 96742 11786
rect 96742 11734 96794 11786
rect 96794 11734 96796 11786
rect 96740 11732 96796 11734
rect 96844 11786 96900 11788
rect 96844 11734 96846 11786
rect 96846 11734 96898 11786
rect 96898 11734 96900 11786
rect 96844 11732 96900 11734
rect 96636 10218 96692 10220
rect 96636 10166 96638 10218
rect 96638 10166 96690 10218
rect 96690 10166 96692 10218
rect 96636 10164 96692 10166
rect 96740 10218 96796 10220
rect 96740 10166 96742 10218
rect 96742 10166 96794 10218
rect 96794 10166 96796 10218
rect 96740 10164 96796 10166
rect 96844 10218 96900 10220
rect 96844 10166 96846 10218
rect 96846 10166 96898 10218
rect 96898 10166 96900 10218
rect 96844 10164 96900 10166
rect 96636 8650 96692 8652
rect 96636 8598 96638 8650
rect 96638 8598 96690 8650
rect 96690 8598 96692 8650
rect 96636 8596 96692 8598
rect 96740 8650 96796 8652
rect 96740 8598 96742 8650
rect 96742 8598 96794 8650
rect 96794 8598 96796 8650
rect 96740 8596 96796 8598
rect 96844 8650 96900 8652
rect 96844 8598 96846 8650
rect 96846 8598 96898 8650
rect 96898 8598 96900 8650
rect 96844 8596 96900 8598
rect 96636 7082 96692 7084
rect 96636 7030 96638 7082
rect 96638 7030 96690 7082
rect 96690 7030 96692 7082
rect 96636 7028 96692 7030
rect 96740 7082 96796 7084
rect 96740 7030 96742 7082
rect 96742 7030 96794 7082
rect 96794 7030 96796 7082
rect 96740 7028 96796 7030
rect 96844 7082 96900 7084
rect 96844 7030 96846 7082
rect 96846 7030 96898 7082
rect 96898 7030 96900 7082
rect 96844 7028 96900 7030
rect 97468 6860 97524 6916
rect 96636 5514 96692 5516
rect 96636 5462 96638 5514
rect 96638 5462 96690 5514
rect 96690 5462 96692 5514
rect 96636 5460 96692 5462
rect 96740 5514 96796 5516
rect 96740 5462 96742 5514
rect 96742 5462 96794 5514
rect 96794 5462 96796 5514
rect 96740 5460 96796 5462
rect 96844 5514 96900 5516
rect 96844 5462 96846 5514
rect 96846 5462 96898 5514
rect 96898 5462 96900 5514
rect 96844 5460 96900 5462
rect 93996 5180 94052 5236
rect 84252 4284 84308 4340
rect 87052 4338 87108 4340
rect 87052 4286 87054 4338
rect 87054 4286 87106 4338
rect 87106 4286 87108 4338
rect 87052 4284 87108 4286
rect 88060 4284 88116 4340
rect 81276 3162 81332 3164
rect 81276 3110 81278 3162
rect 81278 3110 81330 3162
rect 81330 3110 81332 3162
rect 81276 3108 81332 3110
rect 81380 3162 81436 3164
rect 81380 3110 81382 3162
rect 81382 3110 81434 3162
rect 81434 3110 81436 3162
rect 81380 3108 81436 3110
rect 81484 3162 81540 3164
rect 81484 3110 81486 3162
rect 81486 3110 81538 3162
rect 81538 3110 81540 3162
rect 81484 3108 81540 3110
rect 80556 2268 80612 2324
rect 93436 4284 93492 4340
rect 90188 3724 90244 3780
rect 84364 3388 84420 3444
rect 84924 3442 84980 3444
rect 84924 3390 84926 3442
rect 84926 3390 84978 3442
rect 84978 3390 84980 3442
rect 84924 3388 84980 3390
rect 87388 3388 87444 3444
rect 87388 2492 87444 2548
rect 100044 29314 100100 29316
rect 100044 29262 100046 29314
rect 100046 29262 100098 29314
rect 100098 29262 100100 29314
rect 100044 29260 100100 29262
rect 98588 6076 98644 6132
rect 104412 30210 104468 30212
rect 104412 30158 104414 30210
rect 104414 30158 104466 30210
rect 104466 30158 104468 30210
rect 104412 30156 104468 30158
rect 104972 30210 105028 30212
rect 104972 30158 104974 30210
rect 104974 30158 105026 30210
rect 105026 30158 105028 30210
rect 104972 30156 105028 30158
rect 103740 30098 103796 30100
rect 103740 30046 103742 30098
rect 103742 30046 103794 30098
rect 103794 30046 103796 30098
rect 103740 30044 103796 30046
rect 111996 45498 112052 45500
rect 111996 45446 111998 45498
rect 111998 45446 112050 45498
rect 112050 45446 112052 45498
rect 111996 45444 112052 45446
rect 112100 45498 112156 45500
rect 112100 45446 112102 45498
rect 112102 45446 112154 45498
rect 112154 45446 112156 45498
rect 112100 45444 112156 45446
rect 112204 45498 112260 45500
rect 112204 45446 112206 45498
rect 112206 45446 112258 45498
rect 112258 45446 112260 45498
rect 112204 45444 112260 45446
rect 111996 43930 112052 43932
rect 111996 43878 111998 43930
rect 111998 43878 112050 43930
rect 112050 43878 112052 43930
rect 111996 43876 112052 43878
rect 112100 43930 112156 43932
rect 112100 43878 112102 43930
rect 112102 43878 112154 43930
rect 112154 43878 112156 43930
rect 112100 43876 112156 43878
rect 112204 43930 112260 43932
rect 112204 43878 112206 43930
rect 112206 43878 112258 43930
rect 112258 43878 112260 43930
rect 112204 43876 112260 43878
rect 111996 42362 112052 42364
rect 111996 42310 111998 42362
rect 111998 42310 112050 42362
rect 112050 42310 112052 42362
rect 111996 42308 112052 42310
rect 112100 42362 112156 42364
rect 112100 42310 112102 42362
rect 112102 42310 112154 42362
rect 112154 42310 112156 42362
rect 112100 42308 112156 42310
rect 112204 42362 112260 42364
rect 112204 42310 112206 42362
rect 112206 42310 112258 42362
rect 112258 42310 112260 42362
rect 112204 42308 112260 42310
rect 111996 40794 112052 40796
rect 111996 40742 111998 40794
rect 111998 40742 112050 40794
rect 112050 40742 112052 40794
rect 111996 40740 112052 40742
rect 112100 40794 112156 40796
rect 112100 40742 112102 40794
rect 112102 40742 112154 40794
rect 112154 40742 112156 40794
rect 112100 40740 112156 40742
rect 112204 40794 112260 40796
rect 112204 40742 112206 40794
rect 112206 40742 112258 40794
rect 112258 40742 112260 40794
rect 112204 40740 112260 40742
rect 111996 39226 112052 39228
rect 111996 39174 111998 39226
rect 111998 39174 112050 39226
rect 112050 39174 112052 39226
rect 111996 39172 112052 39174
rect 112100 39226 112156 39228
rect 112100 39174 112102 39226
rect 112102 39174 112154 39226
rect 112154 39174 112156 39226
rect 112100 39172 112156 39174
rect 112204 39226 112260 39228
rect 112204 39174 112206 39226
rect 112206 39174 112258 39226
rect 112258 39174 112260 39226
rect 112204 39172 112260 39174
rect 111996 37658 112052 37660
rect 111996 37606 111998 37658
rect 111998 37606 112050 37658
rect 112050 37606 112052 37658
rect 111996 37604 112052 37606
rect 112100 37658 112156 37660
rect 112100 37606 112102 37658
rect 112102 37606 112154 37658
rect 112154 37606 112156 37658
rect 112100 37604 112156 37606
rect 112204 37658 112260 37660
rect 112204 37606 112206 37658
rect 112206 37606 112258 37658
rect 112258 37606 112260 37658
rect 112204 37604 112260 37606
rect 111996 36090 112052 36092
rect 111996 36038 111998 36090
rect 111998 36038 112050 36090
rect 112050 36038 112052 36090
rect 111996 36036 112052 36038
rect 112100 36090 112156 36092
rect 112100 36038 112102 36090
rect 112102 36038 112154 36090
rect 112154 36038 112156 36090
rect 112100 36036 112156 36038
rect 112204 36090 112260 36092
rect 112204 36038 112206 36090
rect 112206 36038 112258 36090
rect 112258 36038 112260 36090
rect 112204 36036 112260 36038
rect 111996 34522 112052 34524
rect 111996 34470 111998 34522
rect 111998 34470 112050 34522
rect 112050 34470 112052 34522
rect 111996 34468 112052 34470
rect 112100 34522 112156 34524
rect 112100 34470 112102 34522
rect 112102 34470 112154 34522
rect 112154 34470 112156 34522
rect 112100 34468 112156 34470
rect 112204 34522 112260 34524
rect 112204 34470 112206 34522
rect 112206 34470 112258 34522
rect 112258 34470 112260 34522
rect 112204 34468 112260 34470
rect 111996 32954 112052 32956
rect 111996 32902 111998 32954
rect 111998 32902 112050 32954
rect 112050 32902 112052 32954
rect 111996 32900 112052 32902
rect 112100 32954 112156 32956
rect 112100 32902 112102 32954
rect 112102 32902 112154 32954
rect 112154 32902 112156 32954
rect 112100 32900 112156 32902
rect 112204 32954 112260 32956
rect 112204 32902 112206 32954
rect 112206 32902 112258 32954
rect 112258 32902 112260 32954
rect 112204 32900 112260 32902
rect 105420 30098 105476 30100
rect 105420 30046 105422 30098
rect 105422 30046 105474 30098
rect 105474 30046 105476 30098
rect 105420 30044 105476 30046
rect 106540 30828 106596 30884
rect 101724 29314 101780 29316
rect 101724 29262 101726 29314
rect 101726 29262 101778 29314
rect 101778 29262 101780 29314
rect 101724 29260 101780 29262
rect 105532 6748 105588 6804
rect 108220 30882 108276 30884
rect 108220 30830 108222 30882
rect 108222 30830 108274 30882
rect 108274 30830 108276 30882
rect 108220 30828 108276 30830
rect 109900 30882 109956 30884
rect 109900 30830 109902 30882
rect 109902 30830 109954 30882
rect 109954 30830 109956 30882
rect 109900 30828 109956 30830
rect 108892 30268 108948 30324
rect 110796 30044 110852 30100
rect 110348 8988 110404 9044
rect 106764 6524 106820 6580
rect 96636 3946 96692 3948
rect 96636 3894 96638 3946
rect 96638 3894 96690 3946
rect 96690 3894 96692 3946
rect 96636 3892 96692 3894
rect 96740 3946 96796 3948
rect 96740 3894 96742 3946
rect 96742 3894 96794 3946
rect 96794 3894 96796 3946
rect 96740 3892 96796 3894
rect 96844 3946 96900 3948
rect 96844 3894 96846 3946
rect 96846 3894 96898 3946
rect 96898 3894 96900 3946
rect 96844 3892 96900 3894
rect 93996 3612 94052 3668
rect 95564 3612 95620 3668
rect 101052 4508 101108 4564
rect 103628 4060 103684 4116
rect 101052 3500 101108 3556
rect 109228 5234 109284 5236
rect 109228 5182 109230 5234
rect 109230 5182 109282 5234
rect 109282 5182 109284 5234
rect 109228 5180 109284 5182
rect 109900 5180 109956 5236
rect 109004 5068 109060 5124
rect 111996 31386 112052 31388
rect 111996 31334 111998 31386
rect 111998 31334 112050 31386
rect 112050 31334 112052 31386
rect 111996 31332 112052 31334
rect 112100 31386 112156 31388
rect 112100 31334 112102 31386
rect 112102 31334 112154 31386
rect 112154 31334 112156 31386
rect 112100 31332 112156 31334
rect 112204 31386 112260 31388
rect 112204 31334 112206 31386
rect 112206 31334 112258 31386
rect 112258 31334 112260 31386
rect 112204 31332 112260 31334
rect 118412 41132 118468 41188
rect 117180 36204 117236 36260
rect 113596 30882 113652 30884
rect 113596 30830 113598 30882
rect 113598 30830 113650 30882
rect 113650 30830 113652 30882
rect 113596 30828 113652 30830
rect 113372 30322 113428 30324
rect 113372 30270 113374 30322
rect 113374 30270 113426 30322
rect 113426 30270 113428 30322
rect 113372 30268 113428 30270
rect 112364 30210 112420 30212
rect 112364 30158 112366 30210
rect 112366 30158 112418 30210
rect 112418 30158 112420 30210
rect 112364 30156 112420 30158
rect 111692 30098 111748 30100
rect 111692 30046 111694 30098
rect 111694 30046 111746 30098
rect 111746 30046 111748 30098
rect 111692 30044 111748 30046
rect 112924 30098 112980 30100
rect 112924 30046 112926 30098
rect 112926 30046 112978 30098
rect 112978 30046 112980 30098
rect 112924 30044 112980 30046
rect 111996 29818 112052 29820
rect 111996 29766 111998 29818
rect 111998 29766 112050 29818
rect 112050 29766 112052 29818
rect 111996 29764 112052 29766
rect 112100 29818 112156 29820
rect 112100 29766 112102 29818
rect 112102 29766 112154 29818
rect 112154 29766 112156 29818
rect 112100 29764 112156 29766
rect 112204 29818 112260 29820
rect 112204 29766 112206 29818
rect 112206 29766 112258 29818
rect 112258 29766 112260 29818
rect 112204 29764 112260 29766
rect 111996 28250 112052 28252
rect 111996 28198 111998 28250
rect 111998 28198 112050 28250
rect 112050 28198 112052 28250
rect 111996 28196 112052 28198
rect 112100 28250 112156 28252
rect 112100 28198 112102 28250
rect 112102 28198 112154 28250
rect 112154 28198 112156 28250
rect 112100 28196 112156 28198
rect 112204 28250 112260 28252
rect 112204 28198 112206 28250
rect 112206 28198 112258 28250
rect 112258 28198 112260 28250
rect 112204 28196 112260 28198
rect 111996 26682 112052 26684
rect 111996 26630 111998 26682
rect 111998 26630 112050 26682
rect 112050 26630 112052 26682
rect 111996 26628 112052 26630
rect 112100 26682 112156 26684
rect 112100 26630 112102 26682
rect 112102 26630 112154 26682
rect 112154 26630 112156 26682
rect 112100 26628 112156 26630
rect 112204 26682 112260 26684
rect 112204 26630 112206 26682
rect 112206 26630 112258 26682
rect 112258 26630 112260 26682
rect 112204 26628 112260 26630
rect 111996 25114 112052 25116
rect 111996 25062 111998 25114
rect 111998 25062 112050 25114
rect 112050 25062 112052 25114
rect 111996 25060 112052 25062
rect 112100 25114 112156 25116
rect 112100 25062 112102 25114
rect 112102 25062 112154 25114
rect 112154 25062 112156 25114
rect 112100 25060 112156 25062
rect 112204 25114 112260 25116
rect 112204 25062 112206 25114
rect 112206 25062 112258 25114
rect 112258 25062 112260 25114
rect 112204 25060 112260 25062
rect 111996 23546 112052 23548
rect 111996 23494 111998 23546
rect 111998 23494 112050 23546
rect 112050 23494 112052 23546
rect 111996 23492 112052 23494
rect 112100 23546 112156 23548
rect 112100 23494 112102 23546
rect 112102 23494 112154 23546
rect 112154 23494 112156 23546
rect 112100 23492 112156 23494
rect 112204 23546 112260 23548
rect 112204 23494 112206 23546
rect 112206 23494 112258 23546
rect 112258 23494 112260 23546
rect 112204 23492 112260 23494
rect 111996 21978 112052 21980
rect 111996 21926 111998 21978
rect 111998 21926 112050 21978
rect 112050 21926 112052 21978
rect 111996 21924 112052 21926
rect 112100 21978 112156 21980
rect 112100 21926 112102 21978
rect 112102 21926 112154 21978
rect 112154 21926 112156 21978
rect 112100 21924 112156 21926
rect 112204 21978 112260 21980
rect 112204 21926 112206 21978
rect 112206 21926 112258 21978
rect 112258 21926 112260 21978
rect 112204 21924 112260 21926
rect 111996 20410 112052 20412
rect 111996 20358 111998 20410
rect 111998 20358 112050 20410
rect 112050 20358 112052 20410
rect 111996 20356 112052 20358
rect 112100 20410 112156 20412
rect 112100 20358 112102 20410
rect 112102 20358 112154 20410
rect 112154 20358 112156 20410
rect 112100 20356 112156 20358
rect 112204 20410 112260 20412
rect 112204 20358 112206 20410
rect 112206 20358 112258 20410
rect 112258 20358 112260 20410
rect 112204 20356 112260 20358
rect 111996 18842 112052 18844
rect 111996 18790 111998 18842
rect 111998 18790 112050 18842
rect 112050 18790 112052 18842
rect 111996 18788 112052 18790
rect 112100 18842 112156 18844
rect 112100 18790 112102 18842
rect 112102 18790 112154 18842
rect 112154 18790 112156 18842
rect 112100 18788 112156 18790
rect 112204 18842 112260 18844
rect 112204 18790 112206 18842
rect 112206 18790 112258 18842
rect 112258 18790 112260 18842
rect 112204 18788 112260 18790
rect 111996 17274 112052 17276
rect 111996 17222 111998 17274
rect 111998 17222 112050 17274
rect 112050 17222 112052 17274
rect 111996 17220 112052 17222
rect 112100 17274 112156 17276
rect 112100 17222 112102 17274
rect 112102 17222 112154 17274
rect 112154 17222 112156 17274
rect 112100 17220 112156 17222
rect 112204 17274 112260 17276
rect 112204 17222 112206 17274
rect 112206 17222 112258 17274
rect 112258 17222 112260 17274
rect 112204 17220 112260 17222
rect 111996 15706 112052 15708
rect 111996 15654 111998 15706
rect 111998 15654 112050 15706
rect 112050 15654 112052 15706
rect 111996 15652 112052 15654
rect 112100 15706 112156 15708
rect 112100 15654 112102 15706
rect 112102 15654 112154 15706
rect 112154 15654 112156 15706
rect 112100 15652 112156 15654
rect 112204 15706 112260 15708
rect 112204 15654 112206 15706
rect 112206 15654 112258 15706
rect 112258 15654 112260 15706
rect 112204 15652 112260 15654
rect 111996 14138 112052 14140
rect 111996 14086 111998 14138
rect 111998 14086 112050 14138
rect 112050 14086 112052 14138
rect 111996 14084 112052 14086
rect 112100 14138 112156 14140
rect 112100 14086 112102 14138
rect 112102 14086 112154 14138
rect 112154 14086 112156 14138
rect 112100 14084 112156 14086
rect 112204 14138 112260 14140
rect 112204 14086 112206 14138
rect 112206 14086 112258 14138
rect 112258 14086 112260 14138
rect 112204 14084 112260 14086
rect 111996 12570 112052 12572
rect 111996 12518 111998 12570
rect 111998 12518 112050 12570
rect 112050 12518 112052 12570
rect 111996 12516 112052 12518
rect 112100 12570 112156 12572
rect 112100 12518 112102 12570
rect 112102 12518 112154 12570
rect 112154 12518 112156 12570
rect 112100 12516 112156 12518
rect 112204 12570 112260 12572
rect 112204 12518 112206 12570
rect 112206 12518 112258 12570
rect 112258 12518 112260 12570
rect 112204 12516 112260 12518
rect 111996 11002 112052 11004
rect 111996 10950 111998 11002
rect 111998 10950 112050 11002
rect 112050 10950 112052 11002
rect 111996 10948 112052 10950
rect 112100 11002 112156 11004
rect 112100 10950 112102 11002
rect 112102 10950 112154 11002
rect 112154 10950 112156 11002
rect 112100 10948 112156 10950
rect 112204 11002 112260 11004
rect 112204 10950 112206 11002
rect 112206 10950 112258 11002
rect 112258 10950 112260 11002
rect 112204 10948 112260 10950
rect 112588 9884 112644 9940
rect 111996 9434 112052 9436
rect 111996 9382 111998 9434
rect 111998 9382 112050 9434
rect 112050 9382 112052 9434
rect 111996 9380 112052 9382
rect 112100 9434 112156 9436
rect 112100 9382 112102 9434
rect 112102 9382 112154 9434
rect 112154 9382 112156 9434
rect 112100 9380 112156 9382
rect 112204 9434 112260 9436
rect 112204 9382 112206 9434
rect 112206 9382 112258 9434
rect 112258 9382 112260 9434
rect 112204 9380 112260 9382
rect 111996 7866 112052 7868
rect 111996 7814 111998 7866
rect 111998 7814 112050 7866
rect 112050 7814 112052 7866
rect 111996 7812 112052 7814
rect 112100 7866 112156 7868
rect 112100 7814 112102 7866
rect 112102 7814 112154 7866
rect 112154 7814 112156 7866
rect 112100 7812 112156 7814
rect 112204 7866 112260 7868
rect 112204 7814 112206 7866
rect 112206 7814 112258 7866
rect 112258 7814 112260 7866
rect 112204 7812 112260 7814
rect 111996 6298 112052 6300
rect 111996 6246 111998 6298
rect 111998 6246 112050 6298
rect 112050 6246 112052 6298
rect 111996 6244 112052 6246
rect 112100 6298 112156 6300
rect 112100 6246 112102 6298
rect 112102 6246 112154 6298
rect 112154 6246 112156 6298
rect 112100 6244 112156 6246
rect 112204 6298 112260 6300
rect 112204 6246 112206 6298
rect 112206 6246 112258 6298
rect 112258 6246 112260 6298
rect 112204 6244 112260 6246
rect 110796 5234 110852 5236
rect 110796 5182 110798 5234
rect 110798 5182 110850 5234
rect 110850 5182 110852 5234
rect 110796 5180 110852 5182
rect 110012 5122 110068 5124
rect 110012 5070 110014 5122
rect 110014 5070 110066 5122
rect 110066 5070 110068 5122
rect 110012 5068 110068 5070
rect 111996 4730 112052 4732
rect 111996 4678 111998 4730
rect 111998 4678 112050 4730
rect 112050 4678 112052 4730
rect 111996 4676 112052 4678
rect 112100 4730 112156 4732
rect 112100 4678 112102 4730
rect 112102 4678 112154 4730
rect 112154 4678 112156 4730
rect 112100 4676 112156 4678
rect 112204 4730 112260 4732
rect 112204 4678 112206 4730
rect 112206 4678 112258 4730
rect 112258 4678 112260 4730
rect 112204 4676 112260 4678
rect 114492 9660 114548 9716
rect 113372 5964 113428 6020
rect 113932 5180 113988 5236
rect 114380 5234 114436 5236
rect 114380 5182 114382 5234
rect 114382 5182 114434 5234
rect 114434 5182 114436 5234
rect 114380 5180 114436 5182
rect 111996 3162 112052 3164
rect 111996 3110 111998 3162
rect 111998 3110 112050 3162
rect 112050 3110 112052 3162
rect 111996 3108 112052 3110
rect 112100 3162 112156 3164
rect 112100 3110 112102 3162
rect 112102 3110 112154 3162
rect 112154 3110 112156 3162
rect 112100 3108 112156 3110
rect 112204 3162 112260 3164
rect 112204 3110 112206 3162
rect 112206 3110 112258 3162
rect 112258 3110 112260 3162
rect 112204 3108 112260 3110
rect 116732 30828 116788 30884
rect 117628 30828 117684 30884
rect 118748 37154 118804 37156
rect 118748 37102 118750 37154
rect 118750 37102 118802 37154
rect 118802 37102 118804 37154
rect 118748 37100 118804 37102
rect 119308 37100 119364 37156
rect 118412 30828 118468 30884
rect 118748 29932 118804 29988
rect 127356 44714 127412 44716
rect 127356 44662 127358 44714
rect 127358 44662 127410 44714
rect 127410 44662 127412 44714
rect 127356 44660 127412 44662
rect 127460 44714 127516 44716
rect 127460 44662 127462 44714
rect 127462 44662 127514 44714
rect 127514 44662 127516 44714
rect 127460 44660 127516 44662
rect 127564 44714 127620 44716
rect 127564 44662 127566 44714
rect 127566 44662 127618 44714
rect 127618 44662 127620 44714
rect 127564 44660 127620 44662
rect 124236 36204 124292 36260
rect 120428 29932 120484 29988
rect 121324 29986 121380 29988
rect 121324 29934 121326 29986
rect 121326 29934 121378 29986
rect 121378 29934 121380 29986
rect 121324 29932 121380 29934
rect 124460 29596 124516 29652
rect 121772 29260 121828 29316
rect 116060 5180 116116 5236
rect 116844 5180 116900 5236
rect 121212 5852 121268 5908
rect 123676 29314 123732 29316
rect 123676 29262 123678 29314
rect 123678 29262 123730 29314
rect 123730 29262 123732 29314
rect 123676 29260 123732 29262
rect 127356 43146 127412 43148
rect 127356 43094 127358 43146
rect 127358 43094 127410 43146
rect 127410 43094 127412 43146
rect 127356 43092 127412 43094
rect 127460 43146 127516 43148
rect 127460 43094 127462 43146
rect 127462 43094 127514 43146
rect 127514 43094 127516 43146
rect 127460 43092 127516 43094
rect 127564 43146 127620 43148
rect 127564 43094 127566 43146
rect 127566 43094 127618 43146
rect 127618 43094 127620 43146
rect 127564 43092 127620 43094
rect 127356 41578 127412 41580
rect 127356 41526 127358 41578
rect 127358 41526 127410 41578
rect 127410 41526 127412 41578
rect 127356 41524 127412 41526
rect 127460 41578 127516 41580
rect 127460 41526 127462 41578
rect 127462 41526 127514 41578
rect 127514 41526 127516 41578
rect 127460 41524 127516 41526
rect 127564 41578 127620 41580
rect 127564 41526 127566 41578
rect 127566 41526 127618 41578
rect 127618 41526 127620 41578
rect 127564 41524 127620 41526
rect 127356 40010 127412 40012
rect 127356 39958 127358 40010
rect 127358 39958 127410 40010
rect 127410 39958 127412 40010
rect 127356 39956 127412 39958
rect 127460 40010 127516 40012
rect 127460 39958 127462 40010
rect 127462 39958 127514 40010
rect 127514 39958 127516 40010
rect 127460 39956 127516 39958
rect 127564 40010 127620 40012
rect 127564 39958 127566 40010
rect 127566 39958 127618 40010
rect 127618 39958 127620 40010
rect 127564 39956 127620 39958
rect 127356 38442 127412 38444
rect 127356 38390 127358 38442
rect 127358 38390 127410 38442
rect 127410 38390 127412 38442
rect 127356 38388 127412 38390
rect 127460 38442 127516 38444
rect 127460 38390 127462 38442
rect 127462 38390 127514 38442
rect 127514 38390 127516 38442
rect 127460 38388 127516 38390
rect 127564 38442 127620 38444
rect 127564 38390 127566 38442
rect 127566 38390 127618 38442
rect 127618 38390 127620 38442
rect 127564 38388 127620 38390
rect 127356 36874 127412 36876
rect 127356 36822 127358 36874
rect 127358 36822 127410 36874
rect 127410 36822 127412 36874
rect 127356 36820 127412 36822
rect 127460 36874 127516 36876
rect 127460 36822 127462 36874
rect 127462 36822 127514 36874
rect 127514 36822 127516 36874
rect 127460 36820 127516 36822
rect 127564 36874 127620 36876
rect 127564 36822 127566 36874
rect 127566 36822 127618 36874
rect 127618 36822 127620 36874
rect 127564 36820 127620 36822
rect 127356 35306 127412 35308
rect 127356 35254 127358 35306
rect 127358 35254 127410 35306
rect 127410 35254 127412 35306
rect 127356 35252 127412 35254
rect 127460 35306 127516 35308
rect 127460 35254 127462 35306
rect 127462 35254 127514 35306
rect 127514 35254 127516 35306
rect 127460 35252 127516 35254
rect 127564 35306 127620 35308
rect 127564 35254 127566 35306
rect 127566 35254 127618 35306
rect 127618 35254 127620 35306
rect 127564 35252 127620 35254
rect 127356 33738 127412 33740
rect 127356 33686 127358 33738
rect 127358 33686 127410 33738
rect 127410 33686 127412 33738
rect 127356 33684 127412 33686
rect 127460 33738 127516 33740
rect 127460 33686 127462 33738
rect 127462 33686 127514 33738
rect 127514 33686 127516 33738
rect 127460 33684 127516 33686
rect 127564 33738 127620 33740
rect 127564 33686 127566 33738
rect 127566 33686 127618 33738
rect 127618 33686 127620 33738
rect 127564 33684 127620 33686
rect 127356 32170 127412 32172
rect 127356 32118 127358 32170
rect 127358 32118 127410 32170
rect 127410 32118 127412 32170
rect 127356 32116 127412 32118
rect 127460 32170 127516 32172
rect 127460 32118 127462 32170
rect 127462 32118 127514 32170
rect 127514 32118 127516 32170
rect 127460 32116 127516 32118
rect 127564 32170 127620 32172
rect 127564 32118 127566 32170
rect 127566 32118 127618 32170
rect 127618 32118 127620 32170
rect 127564 32116 127620 32118
rect 127356 30602 127412 30604
rect 127356 30550 127358 30602
rect 127358 30550 127410 30602
rect 127410 30550 127412 30602
rect 127356 30548 127412 30550
rect 127460 30602 127516 30604
rect 127460 30550 127462 30602
rect 127462 30550 127514 30602
rect 127514 30550 127516 30602
rect 127460 30548 127516 30550
rect 127564 30602 127620 30604
rect 127564 30550 127566 30602
rect 127566 30550 127618 30602
rect 127618 30550 127620 30602
rect 127564 30548 127620 30550
rect 125356 30156 125412 30212
rect 125356 29650 125412 29652
rect 125356 29598 125358 29650
rect 125358 29598 125410 29650
rect 125410 29598 125412 29650
rect 125356 29596 125412 29598
rect 126140 30044 126196 30100
rect 124908 29314 124964 29316
rect 124908 29262 124910 29314
rect 124910 29262 124962 29314
rect 124962 29262 124964 29314
rect 124908 29260 124964 29262
rect 125580 6412 125636 6468
rect 125132 5964 125188 6020
rect 117628 4844 117684 4900
rect 120092 4172 120148 4228
rect 116844 3724 116900 3780
rect 117068 3724 117124 3780
rect 122444 2380 122500 2436
rect 128940 30210 128996 30212
rect 128940 30158 128942 30210
rect 128942 30158 128994 30210
rect 128994 30158 128996 30210
rect 128940 30156 128996 30158
rect 129948 30210 130004 30212
rect 129948 30158 129950 30210
rect 129950 30158 130002 30210
rect 130002 30158 130004 30210
rect 129948 30156 130004 30158
rect 128268 30098 128324 30100
rect 128268 30046 128270 30098
rect 128270 30046 128322 30098
rect 128322 30046 128324 30098
rect 128268 30044 128324 30046
rect 129500 30098 129556 30100
rect 129500 30046 129502 30098
rect 129502 30046 129554 30098
rect 129554 30046 129556 30098
rect 129500 30044 129556 30046
rect 127356 29034 127412 29036
rect 127356 28982 127358 29034
rect 127358 28982 127410 29034
rect 127410 28982 127412 29034
rect 127356 28980 127412 28982
rect 127460 29034 127516 29036
rect 127460 28982 127462 29034
rect 127462 28982 127514 29034
rect 127514 28982 127516 29034
rect 127460 28980 127516 28982
rect 127564 29034 127620 29036
rect 127564 28982 127566 29034
rect 127566 28982 127618 29034
rect 127618 28982 127620 29034
rect 127564 28980 127620 28982
rect 127356 27466 127412 27468
rect 127356 27414 127358 27466
rect 127358 27414 127410 27466
rect 127410 27414 127412 27466
rect 127356 27412 127412 27414
rect 127460 27466 127516 27468
rect 127460 27414 127462 27466
rect 127462 27414 127514 27466
rect 127514 27414 127516 27466
rect 127460 27412 127516 27414
rect 127564 27466 127620 27468
rect 127564 27414 127566 27466
rect 127566 27414 127618 27466
rect 127618 27414 127620 27466
rect 127564 27412 127620 27414
rect 127356 25898 127412 25900
rect 127356 25846 127358 25898
rect 127358 25846 127410 25898
rect 127410 25846 127412 25898
rect 127356 25844 127412 25846
rect 127460 25898 127516 25900
rect 127460 25846 127462 25898
rect 127462 25846 127514 25898
rect 127514 25846 127516 25898
rect 127460 25844 127516 25846
rect 127564 25898 127620 25900
rect 127564 25846 127566 25898
rect 127566 25846 127618 25898
rect 127618 25846 127620 25898
rect 127564 25844 127620 25846
rect 127356 24330 127412 24332
rect 127356 24278 127358 24330
rect 127358 24278 127410 24330
rect 127410 24278 127412 24330
rect 127356 24276 127412 24278
rect 127460 24330 127516 24332
rect 127460 24278 127462 24330
rect 127462 24278 127514 24330
rect 127514 24278 127516 24330
rect 127460 24276 127516 24278
rect 127564 24330 127620 24332
rect 127564 24278 127566 24330
rect 127566 24278 127618 24330
rect 127618 24278 127620 24330
rect 127564 24276 127620 24278
rect 127356 22762 127412 22764
rect 127356 22710 127358 22762
rect 127358 22710 127410 22762
rect 127410 22710 127412 22762
rect 127356 22708 127412 22710
rect 127460 22762 127516 22764
rect 127460 22710 127462 22762
rect 127462 22710 127514 22762
rect 127514 22710 127516 22762
rect 127460 22708 127516 22710
rect 127564 22762 127620 22764
rect 127564 22710 127566 22762
rect 127566 22710 127618 22762
rect 127618 22710 127620 22762
rect 127564 22708 127620 22710
rect 127356 21194 127412 21196
rect 127356 21142 127358 21194
rect 127358 21142 127410 21194
rect 127410 21142 127412 21194
rect 127356 21140 127412 21142
rect 127460 21194 127516 21196
rect 127460 21142 127462 21194
rect 127462 21142 127514 21194
rect 127514 21142 127516 21194
rect 127460 21140 127516 21142
rect 127564 21194 127620 21196
rect 127564 21142 127566 21194
rect 127566 21142 127618 21194
rect 127618 21142 127620 21194
rect 127564 21140 127620 21142
rect 127356 19626 127412 19628
rect 127356 19574 127358 19626
rect 127358 19574 127410 19626
rect 127410 19574 127412 19626
rect 127356 19572 127412 19574
rect 127460 19626 127516 19628
rect 127460 19574 127462 19626
rect 127462 19574 127514 19626
rect 127514 19574 127516 19626
rect 127460 19572 127516 19574
rect 127564 19626 127620 19628
rect 127564 19574 127566 19626
rect 127566 19574 127618 19626
rect 127618 19574 127620 19626
rect 127564 19572 127620 19574
rect 127356 18058 127412 18060
rect 127356 18006 127358 18058
rect 127358 18006 127410 18058
rect 127410 18006 127412 18058
rect 127356 18004 127412 18006
rect 127460 18058 127516 18060
rect 127460 18006 127462 18058
rect 127462 18006 127514 18058
rect 127514 18006 127516 18058
rect 127460 18004 127516 18006
rect 127564 18058 127620 18060
rect 127564 18006 127566 18058
rect 127566 18006 127618 18058
rect 127618 18006 127620 18058
rect 127564 18004 127620 18006
rect 127356 16490 127412 16492
rect 127356 16438 127358 16490
rect 127358 16438 127410 16490
rect 127410 16438 127412 16490
rect 127356 16436 127412 16438
rect 127460 16490 127516 16492
rect 127460 16438 127462 16490
rect 127462 16438 127514 16490
rect 127514 16438 127516 16490
rect 127460 16436 127516 16438
rect 127564 16490 127620 16492
rect 127564 16438 127566 16490
rect 127566 16438 127618 16490
rect 127618 16438 127620 16490
rect 127564 16436 127620 16438
rect 127356 14922 127412 14924
rect 127356 14870 127358 14922
rect 127358 14870 127410 14922
rect 127410 14870 127412 14922
rect 127356 14868 127412 14870
rect 127460 14922 127516 14924
rect 127460 14870 127462 14922
rect 127462 14870 127514 14922
rect 127514 14870 127516 14922
rect 127460 14868 127516 14870
rect 127564 14922 127620 14924
rect 127564 14870 127566 14922
rect 127566 14870 127618 14922
rect 127618 14870 127620 14922
rect 127564 14868 127620 14870
rect 127356 13354 127412 13356
rect 127356 13302 127358 13354
rect 127358 13302 127410 13354
rect 127410 13302 127412 13354
rect 127356 13300 127412 13302
rect 127460 13354 127516 13356
rect 127460 13302 127462 13354
rect 127462 13302 127514 13354
rect 127514 13302 127516 13354
rect 127460 13300 127516 13302
rect 127564 13354 127620 13356
rect 127564 13302 127566 13354
rect 127566 13302 127618 13354
rect 127618 13302 127620 13354
rect 127564 13300 127620 13302
rect 127356 11786 127412 11788
rect 127356 11734 127358 11786
rect 127358 11734 127410 11786
rect 127410 11734 127412 11786
rect 127356 11732 127412 11734
rect 127460 11786 127516 11788
rect 127460 11734 127462 11786
rect 127462 11734 127514 11786
rect 127514 11734 127516 11786
rect 127460 11732 127516 11734
rect 127564 11786 127620 11788
rect 127564 11734 127566 11786
rect 127566 11734 127618 11786
rect 127618 11734 127620 11786
rect 127564 11732 127620 11734
rect 127356 10218 127412 10220
rect 127356 10166 127358 10218
rect 127358 10166 127410 10218
rect 127410 10166 127412 10218
rect 127356 10164 127412 10166
rect 127460 10218 127516 10220
rect 127460 10166 127462 10218
rect 127462 10166 127514 10218
rect 127514 10166 127516 10218
rect 127460 10164 127516 10166
rect 127564 10218 127620 10220
rect 127564 10166 127566 10218
rect 127566 10166 127618 10218
rect 127618 10166 127620 10218
rect 127564 10164 127620 10166
rect 127356 8650 127412 8652
rect 127356 8598 127358 8650
rect 127358 8598 127410 8650
rect 127410 8598 127412 8650
rect 127356 8596 127412 8598
rect 127460 8650 127516 8652
rect 127460 8598 127462 8650
rect 127462 8598 127514 8650
rect 127514 8598 127516 8650
rect 127460 8596 127516 8598
rect 127564 8650 127620 8652
rect 127564 8598 127566 8650
rect 127566 8598 127618 8650
rect 127618 8598 127620 8650
rect 127564 8596 127620 8598
rect 139916 45612 139972 45668
rect 135660 45164 135716 45220
rect 131964 44322 132020 44324
rect 131964 44270 131966 44322
rect 131966 44270 132018 44322
rect 132018 44270 132020 44322
rect 131964 44268 132020 44270
rect 135100 44322 135156 44324
rect 135100 44270 135102 44322
rect 135102 44270 135154 44322
rect 135154 44270 135156 44322
rect 135100 44268 135156 44270
rect 138124 44994 138180 44996
rect 138124 44942 138126 44994
rect 138126 44942 138178 44994
rect 138178 44942 138180 44994
rect 138124 44940 138180 44942
rect 135772 43538 135828 43540
rect 135772 43486 135774 43538
rect 135774 43486 135826 43538
rect 135826 43486 135828 43538
rect 135772 43484 135828 43486
rect 136108 43484 136164 43540
rect 135100 43426 135156 43428
rect 135100 43374 135102 43426
rect 135102 43374 135154 43426
rect 135154 43374 135156 43426
rect 135100 43372 135156 43374
rect 135996 43372 136052 43428
rect 134764 42700 134820 42756
rect 133980 39452 134036 39508
rect 130508 36258 130564 36260
rect 130508 36206 130510 36258
rect 130510 36206 130562 36258
rect 130562 36206 130564 36258
rect 130508 36204 130564 36206
rect 131068 36204 131124 36260
rect 132636 34636 132692 34692
rect 132860 30210 132916 30212
rect 132860 30158 132862 30210
rect 132862 30158 132914 30210
rect 132914 30158 132916 30210
rect 132860 30156 132916 30158
rect 132636 30044 132692 30100
rect 133644 30098 133700 30100
rect 133644 30046 133646 30098
rect 133646 30046 133698 30098
rect 133698 30046 133700 30098
rect 133644 30044 133700 30046
rect 137228 43426 137284 43428
rect 137228 43374 137230 43426
rect 137230 43374 137282 43426
rect 137282 43374 137284 43426
rect 137228 43372 137284 43374
rect 137564 42924 137620 42980
rect 138684 43484 138740 43540
rect 138124 42978 138180 42980
rect 138124 42926 138126 42978
rect 138126 42926 138178 42978
rect 138178 42926 138180 42978
rect 138124 42924 138180 42926
rect 137900 42754 137956 42756
rect 137900 42702 137902 42754
rect 137902 42702 137954 42754
rect 137954 42702 137956 42754
rect 137900 42700 137956 42702
rect 136220 42476 136276 42532
rect 137788 42530 137844 42532
rect 137788 42478 137790 42530
rect 137790 42478 137842 42530
rect 137842 42478 137844 42530
rect 137788 42476 137844 42478
rect 136108 35196 136164 35252
rect 136780 35196 136836 35252
rect 136332 30882 136388 30884
rect 136332 30830 136334 30882
rect 136334 30830 136386 30882
rect 136386 30830 136388 30882
rect 136332 30828 136388 30830
rect 138124 30882 138180 30884
rect 138124 30830 138126 30882
rect 138126 30830 138178 30882
rect 138178 30830 138180 30882
rect 138124 30828 138180 30830
rect 133980 29650 134036 29652
rect 133980 29598 133982 29650
rect 133982 29598 134034 29650
rect 134034 29598 134036 29650
rect 133980 29596 134036 29598
rect 134428 30156 134484 30212
rect 135772 29596 135828 29652
rect 134652 17612 134708 17668
rect 132748 15932 132804 15988
rect 131068 11228 131124 11284
rect 131068 9100 131124 9156
rect 130172 8316 130228 8372
rect 134540 9042 134596 9044
rect 134540 8990 134542 9042
rect 134542 8990 134594 9042
rect 134594 8990 134596 9042
rect 134540 8988 134596 8990
rect 132860 8370 132916 8372
rect 132860 8318 132862 8370
rect 132862 8318 132914 8370
rect 132914 8318 132916 8370
rect 132860 8316 132916 8318
rect 132524 7586 132580 7588
rect 132524 7534 132526 7586
rect 132526 7534 132578 7586
rect 132578 7534 132580 7586
rect 132524 7532 132580 7534
rect 130508 7420 130564 7476
rect 127356 7082 127412 7084
rect 127356 7030 127358 7082
rect 127358 7030 127410 7082
rect 127410 7030 127412 7082
rect 127356 7028 127412 7030
rect 127460 7082 127516 7084
rect 127460 7030 127462 7082
rect 127462 7030 127514 7082
rect 127514 7030 127516 7082
rect 127460 7028 127516 7030
rect 127564 7082 127620 7084
rect 127564 7030 127566 7082
rect 127566 7030 127618 7082
rect 127618 7030 127620 7082
rect 127564 7028 127620 7030
rect 130060 6076 130116 6132
rect 127356 5514 127412 5516
rect 127356 5462 127358 5514
rect 127358 5462 127410 5514
rect 127410 5462 127412 5514
rect 127356 5460 127412 5462
rect 127460 5514 127516 5516
rect 127460 5462 127462 5514
rect 127462 5462 127514 5514
rect 127514 5462 127516 5514
rect 127460 5460 127516 5462
rect 127564 5514 127620 5516
rect 127564 5462 127566 5514
rect 127566 5462 127618 5514
rect 127618 5462 127620 5514
rect 127564 5460 127620 5462
rect 131740 7474 131796 7476
rect 131740 7422 131742 7474
rect 131742 7422 131794 7474
rect 131794 7422 131796 7474
rect 131740 7420 131796 7422
rect 131964 7420 132020 7476
rect 131740 6860 131796 6916
rect 131292 6636 131348 6692
rect 127820 4620 127876 4676
rect 127356 3946 127412 3948
rect 127356 3894 127358 3946
rect 127358 3894 127410 3946
rect 127410 3894 127412 3946
rect 127356 3892 127412 3894
rect 127460 3946 127516 3948
rect 127460 3894 127462 3946
rect 127462 3894 127514 3946
rect 127514 3894 127516 3946
rect 127460 3892 127516 3894
rect 127564 3946 127620 3948
rect 127564 3894 127566 3946
rect 127566 3894 127618 3946
rect 127618 3894 127620 3946
rect 127564 3892 127620 3894
rect 130508 4508 130564 4564
rect 134316 8204 134372 8260
rect 133084 6860 133140 6916
rect 133196 7532 133252 7588
rect 133084 6690 133140 6692
rect 133084 6638 133086 6690
rect 133086 6638 133138 6690
rect 133138 6638 133140 6690
rect 133084 6636 133140 6638
rect 132076 6524 132132 6580
rect 133756 6076 133812 6132
rect 134204 6860 134260 6916
rect 133980 5852 134036 5908
rect 134540 7532 134596 7588
rect 136220 30210 136276 30212
rect 136220 30158 136222 30210
rect 136222 30158 136274 30210
rect 136274 30158 136276 30210
rect 136220 30156 136276 30158
rect 136780 30156 136836 30212
rect 135884 10444 135940 10500
rect 136220 19292 136276 19348
rect 135324 9154 135380 9156
rect 135324 9102 135326 9154
rect 135326 9102 135378 9154
rect 135378 9102 135380 9154
rect 135324 9100 135380 9102
rect 135996 9154 136052 9156
rect 135996 9102 135998 9154
rect 135998 9102 136050 9154
rect 136050 9102 136052 9154
rect 135996 9100 136052 9102
rect 135548 9042 135604 9044
rect 135548 8990 135550 9042
rect 135550 8990 135602 9042
rect 135602 8990 135604 9042
rect 135548 8988 135604 8990
rect 135772 8146 135828 8148
rect 135772 8094 135774 8146
rect 135774 8094 135826 8146
rect 135826 8094 135828 8146
rect 135772 8092 135828 8094
rect 135548 7980 135604 8036
rect 139804 44994 139860 44996
rect 139804 44942 139806 44994
rect 139806 44942 139858 44994
rect 139858 44942 139860 44994
rect 139804 44940 139860 44942
rect 144284 45666 144340 45668
rect 144284 45614 144286 45666
rect 144286 45614 144338 45666
rect 144338 45614 144340 45666
rect 144284 45612 144340 45614
rect 142716 45498 142772 45500
rect 142716 45446 142718 45498
rect 142718 45446 142770 45498
rect 142770 45446 142772 45498
rect 142716 45444 142772 45446
rect 142820 45498 142876 45500
rect 142820 45446 142822 45498
rect 142822 45446 142874 45498
rect 142874 45446 142876 45498
rect 142820 45444 142876 45446
rect 142924 45498 142980 45500
rect 142924 45446 142926 45498
rect 142926 45446 142978 45498
rect 142978 45446 142980 45498
rect 142924 45444 142980 45446
rect 140588 45218 140644 45220
rect 140588 45166 140590 45218
rect 140590 45166 140642 45218
rect 140642 45166 140644 45218
rect 140588 45164 140644 45166
rect 141932 44940 141988 44996
rect 140364 43538 140420 43540
rect 140364 43486 140366 43538
rect 140366 43486 140418 43538
rect 140418 43486 140420 43538
rect 140364 43484 140420 43486
rect 137900 11452 137956 11508
rect 138012 14252 138068 14308
rect 137676 10332 137732 10388
rect 136332 8092 136388 8148
rect 135660 7586 135716 7588
rect 135660 7534 135662 7586
rect 135662 7534 135714 7586
rect 135714 7534 135716 7586
rect 135660 7532 135716 7534
rect 135548 7474 135604 7476
rect 135548 7422 135550 7474
rect 135550 7422 135602 7474
rect 135602 7422 135604 7474
rect 135548 7420 135604 7422
rect 135100 5852 135156 5908
rect 133420 5234 133476 5236
rect 133420 5182 133422 5234
rect 133422 5182 133474 5234
rect 133474 5182 133476 5234
rect 133420 5180 133476 5182
rect 132972 4284 133028 4340
rect 130844 4060 130900 4116
rect 132972 4060 133028 4116
rect 133196 4284 133252 4340
rect 131292 3500 131348 3556
rect 133756 4060 133812 4116
rect 135548 6636 135604 6692
rect 136332 6690 136388 6692
rect 136332 6638 136334 6690
rect 136334 6638 136386 6690
rect 136386 6638 136388 6690
rect 136332 6636 136388 6638
rect 135772 6412 135828 6468
rect 135772 5346 135828 5348
rect 135772 5294 135774 5346
rect 135774 5294 135826 5346
rect 135826 5294 135828 5346
rect 135772 5292 135828 5294
rect 136444 5292 136500 5348
rect 135324 4732 135380 4788
rect 135884 4956 135940 5012
rect 135324 3612 135380 3668
rect 135100 2940 135156 2996
rect 136444 4396 136500 4452
rect 137676 7532 137732 7588
rect 137228 6748 137284 6804
rect 137900 6466 137956 6468
rect 137900 6414 137902 6466
rect 137902 6414 137954 6466
rect 137954 6414 137956 6466
rect 137900 6412 137956 6414
rect 139132 11564 139188 11620
rect 138460 10780 138516 10836
rect 138236 10108 138292 10164
rect 138124 9100 138180 9156
rect 139132 10108 139188 10164
rect 138684 9996 138740 10052
rect 140252 13468 140308 13524
rect 140140 12684 140196 12740
rect 140028 11116 140084 11172
rect 138684 9100 138740 9156
rect 139132 9100 139188 9156
rect 139804 9100 139860 9156
rect 139468 8258 139524 8260
rect 139468 8206 139470 8258
rect 139470 8206 139522 8258
rect 139522 8206 139524 8258
rect 139468 8204 139524 8206
rect 138236 6690 138292 6692
rect 138236 6638 138238 6690
rect 138238 6638 138290 6690
rect 138290 6638 138292 6690
rect 138236 6636 138292 6638
rect 137452 5234 137508 5236
rect 137452 5182 137454 5234
rect 137454 5182 137506 5234
rect 137506 5182 137508 5234
rect 137452 5180 137508 5182
rect 138124 5122 138180 5124
rect 138124 5070 138126 5122
rect 138126 5070 138178 5122
rect 138178 5070 138180 5122
rect 138124 5068 138180 5070
rect 137004 4844 137060 4900
rect 138908 4956 138964 5012
rect 139132 6076 139188 6132
rect 139244 7420 139300 7476
rect 139132 5906 139188 5908
rect 139132 5854 139134 5906
rect 139134 5854 139186 5906
rect 139186 5854 139188 5906
rect 139132 5852 139188 5854
rect 138012 4844 138068 4900
rect 138796 4844 138852 4900
rect 138124 4620 138180 4676
rect 137340 4338 137396 4340
rect 137340 4286 137342 4338
rect 137342 4286 137394 4338
rect 137394 4286 137396 4338
rect 137340 4284 137396 4286
rect 136556 2716 136612 2772
rect 139468 6748 139524 6804
rect 139356 6412 139412 6468
rect 140924 9212 140980 9268
rect 140252 9154 140308 9156
rect 140252 9102 140254 9154
rect 140254 9102 140306 9154
rect 140306 9102 140308 9154
rect 140252 9100 140308 9102
rect 140812 7644 140868 7700
rect 140588 7474 140644 7476
rect 140588 7422 140590 7474
rect 140590 7422 140642 7474
rect 140642 7422 140644 7474
rect 140588 7420 140644 7422
rect 139468 5794 139524 5796
rect 139468 5742 139470 5794
rect 139470 5742 139522 5794
rect 139522 5742 139524 5794
rect 139468 5740 139524 5742
rect 140364 6578 140420 6580
rect 140364 6526 140366 6578
rect 140366 6526 140418 6578
rect 140418 6526 140420 6578
rect 140364 6524 140420 6526
rect 140588 5794 140644 5796
rect 140588 5742 140590 5794
rect 140590 5742 140642 5794
rect 140642 5742 140644 5794
rect 140588 5740 140644 5742
rect 140364 4844 140420 4900
rect 140476 5068 140532 5124
rect 139804 4620 139860 4676
rect 141036 5740 141092 5796
rect 140252 4172 140308 4228
rect 140924 3612 140980 3668
rect 139356 2828 139412 2884
rect 141260 5068 141316 5124
rect 142716 43930 142772 43932
rect 142716 43878 142718 43930
rect 142718 43878 142770 43930
rect 142770 43878 142772 43930
rect 142716 43876 142772 43878
rect 142820 43930 142876 43932
rect 142820 43878 142822 43930
rect 142822 43878 142874 43930
rect 142874 43878 142876 43930
rect 142820 43876 142876 43878
rect 142924 43930 142980 43932
rect 142924 43878 142926 43930
rect 142926 43878 142978 43930
rect 142978 43878 142980 43930
rect 142924 43876 142980 43878
rect 142716 42362 142772 42364
rect 142716 42310 142718 42362
rect 142718 42310 142770 42362
rect 142770 42310 142772 42362
rect 142716 42308 142772 42310
rect 142820 42362 142876 42364
rect 142820 42310 142822 42362
rect 142822 42310 142874 42362
rect 142874 42310 142876 42362
rect 142820 42308 142876 42310
rect 142924 42362 142980 42364
rect 142924 42310 142926 42362
rect 142926 42310 142978 42362
rect 142978 42310 142980 42362
rect 142924 42308 142980 42310
rect 142716 40794 142772 40796
rect 142716 40742 142718 40794
rect 142718 40742 142770 40794
rect 142770 40742 142772 40794
rect 142716 40740 142772 40742
rect 142820 40794 142876 40796
rect 142820 40742 142822 40794
rect 142822 40742 142874 40794
rect 142874 40742 142876 40794
rect 142820 40740 142876 40742
rect 142924 40794 142980 40796
rect 142924 40742 142926 40794
rect 142926 40742 142978 40794
rect 142978 40742 142980 40794
rect 142924 40740 142980 40742
rect 142716 39226 142772 39228
rect 142716 39174 142718 39226
rect 142718 39174 142770 39226
rect 142770 39174 142772 39226
rect 142716 39172 142772 39174
rect 142820 39226 142876 39228
rect 142820 39174 142822 39226
rect 142822 39174 142874 39226
rect 142874 39174 142876 39226
rect 142820 39172 142876 39174
rect 142924 39226 142980 39228
rect 142924 39174 142926 39226
rect 142926 39174 142978 39226
rect 142978 39174 142980 39226
rect 142924 39172 142980 39174
rect 142716 37658 142772 37660
rect 142716 37606 142718 37658
rect 142718 37606 142770 37658
rect 142770 37606 142772 37658
rect 142716 37604 142772 37606
rect 142820 37658 142876 37660
rect 142820 37606 142822 37658
rect 142822 37606 142874 37658
rect 142874 37606 142876 37658
rect 142820 37604 142876 37606
rect 142924 37658 142980 37660
rect 142924 37606 142926 37658
rect 142926 37606 142978 37658
rect 142978 37606 142980 37658
rect 142924 37604 142980 37606
rect 142716 36090 142772 36092
rect 142716 36038 142718 36090
rect 142718 36038 142770 36090
rect 142770 36038 142772 36090
rect 142716 36036 142772 36038
rect 142820 36090 142876 36092
rect 142820 36038 142822 36090
rect 142822 36038 142874 36090
rect 142874 36038 142876 36090
rect 142820 36036 142876 36038
rect 142924 36090 142980 36092
rect 142924 36038 142926 36090
rect 142926 36038 142978 36090
rect 142978 36038 142980 36090
rect 142924 36036 142980 36038
rect 142716 34522 142772 34524
rect 142716 34470 142718 34522
rect 142718 34470 142770 34522
rect 142770 34470 142772 34522
rect 142716 34468 142772 34470
rect 142820 34522 142876 34524
rect 142820 34470 142822 34522
rect 142822 34470 142874 34522
rect 142874 34470 142876 34522
rect 142820 34468 142876 34470
rect 142924 34522 142980 34524
rect 142924 34470 142926 34522
rect 142926 34470 142978 34522
rect 142978 34470 142980 34522
rect 142924 34468 142980 34470
rect 142716 32954 142772 32956
rect 142716 32902 142718 32954
rect 142718 32902 142770 32954
rect 142770 32902 142772 32954
rect 142716 32900 142772 32902
rect 142820 32954 142876 32956
rect 142820 32902 142822 32954
rect 142822 32902 142874 32954
rect 142874 32902 142876 32954
rect 142820 32900 142876 32902
rect 142924 32954 142980 32956
rect 142924 32902 142926 32954
rect 142926 32902 142978 32954
rect 142978 32902 142980 32954
rect 142924 32900 142980 32902
rect 142716 31386 142772 31388
rect 142716 31334 142718 31386
rect 142718 31334 142770 31386
rect 142770 31334 142772 31386
rect 142716 31332 142772 31334
rect 142820 31386 142876 31388
rect 142820 31334 142822 31386
rect 142822 31334 142874 31386
rect 142874 31334 142876 31386
rect 142820 31332 142876 31334
rect 142924 31386 142980 31388
rect 142924 31334 142926 31386
rect 142926 31334 142978 31386
rect 142978 31334 142980 31386
rect 142924 31332 142980 31334
rect 142716 29818 142772 29820
rect 142716 29766 142718 29818
rect 142718 29766 142770 29818
rect 142770 29766 142772 29818
rect 142716 29764 142772 29766
rect 142820 29818 142876 29820
rect 142820 29766 142822 29818
rect 142822 29766 142874 29818
rect 142874 29766 142876 29818
rect 142820 29764 142876 29766
rect 142924 29818 142980 29820
rect 142924 29766 142926 29818
rect 142926 29766 142978 29818
rect 142978 29766 142980 29818
rect 142924 29764 142980 29766
rect 142716 28250 142772 28252
rect 142716 28198 142718 28250
rect 142718 28198 142770 28250
rect 142770 28198 142772 28250
rect 142716 28196 142772 28198
rect 142820 28250 142876 28252
rect 142820 28198 142822 28250
rect 142822 28198 142874 28250
rect 142874 28198 142876 28250
rect 142820 28196 142876 28198
rect 142924 28250 142980 28252
rect 142924 28198 142926 28250
rect 142926 28198 142978 28250
rect 142978 28198 142980 28250
rect 142924 28196 142980 28198
rect 142716 26682 142772 26684
rect 142716 26630 142718 26682
rect 142718 26630 142770 26682
rect 142770 26630 142772 26682
rect 142716 26628 142772 26630
rect 142820 26682 142876 26684
rect 142820 26630 142822 26682
rect 142822 26630 142874 26682
rect 142874 26630 142876 26682
rect 142820 26628 142876 26630
rect 142924 26682 142980 26684
rect 142924 26630 142926 26682
rect 142926 26630 142978 26682
rect 142978 26630 142980 26682
rect 142924 26628 142980 26630
rect 142716 25114 142772 25116
rect 142716 25062 142718 25114
rect 142718 25062 142770 25114
rect 142770 25062 142772 25114
rect 142716 25060 142772 25062
rect 142820 25114 142876 25116
rect 142820 25062 142822 25114
rect 142822 25062 142874 25114
rect 142874 25062 142876 25114
rect 142820 25060 142876 25062
rect 142924 25114 142980 25116
rect 142924 25062 142926 25114
rect 142926 25062 142978 25114
rect 142978 25062 142980 25114
rect 142924 25060 142980 25062
rect 142716 23546 142772 23548
rect 142716 23494 142718 23546
rect 142718 23494 142770 23546
rect 142770 23494 142772 23546
rect 142716 23492 142772 23494
rect 142820 23546 142876 23548
rect 142820 23494 142822 23546
rect 142822 23494 142874 23546
rect 142874 23494 142876 23546
rect 142820 23492 142876 23494
rect 142924 23546 142980 23548
rect 142924 23494 142926 23546
rect 142926 23494 142978 23546
rect 142978 23494 142980 23546
rect 142924 23492 142980 23494
rect 142716 21978 142772 21980
rect 142716 21926 142718 21978
rect 142718 21926 142770 21978
rect 142770 21926 142772 21978
rect 142716 21924 142772 21926
rect 142820 21978 142876 21980
rect 142820 21926 142822 21978
rect 142822 21926 142874 21978
rect 142874 21926 142876 21978
rect 142820 21924 142876 21926
rect 142924 21978 142980 21980
rect 142924 21926 142926 21978
rect 142926 21926 142978 21978
rect 142978 21926 142980 21978
rect 142924 21924 142980 21926
rect 142716 20410 142772 20412
rect 142716 20358 142718 20410
rect 142718 20358 142770 20410
rect 142770 20358 142772 20410
rect 142716 20356 142772 20358
rect 142820 20410 142876 20412
rect 142820 20358 142822 20410
rect 142822 20358 142874 20410
rect 142874 20358 142876 20410
rect 142820 20356 142876 20358
rect 142924 20410 142980 20412
rect 142924 20358 142926 20410
rect 142926 20358 142978 20410
rect 142978 20358 142980 20410
rect 142924 20356 142980 20358
rect 142716 18842 142772 18844
rect 142716 18790 142718 18842
rect 142718 18790 142770 18842
rect 142770 18790 142772 18842
rect 142716 18788 142772 18790
rect 142820 18842 142876 18844
rect 142820 18790 142822 18842
rect 142822 18790 142874 18842
rect 142874 18790 142876 18842
rect 142820 18788 142876 18790
rect 142924 18842 142980 18844
rect 142924 18790 142926 18842
rect 142926 18790 142978 18842
rect 142978 18790 142980 18842
rect 142924 18788 142980 18790
rect 145852 17612 145908 17668
rect 142716 17274 142772 17276
rect 142716 17222 142718 17274
rect 142718 17222 142770 17274
rect 142770 17222 142772 17274
rect 142716 17220 142772 17222
rect 142820 17274 142876 17276
rect 142820 17222 142822 17274
rect 142822 17222 142874 17274
rect 142874 17222 142876 17274
rect 142820 17220 142876 17222
rect 142924 17274 142980 17276
rect 142924 17222 142926 17274
rect 142926 17222 142978 17274
rect 142978 17222 142980 17274
rect 142924 17220 142980 17222
rect 142716 15706 142772 15708
rect 142716 15654 142718 15706
rect 142718 15654 142770 15706
rect 142770 15654 142772 15706
rect 142716 15652 142772 15654
rect 142820 15706 142876 15708
rect 142820 15654 142822 15706
rect 142822 15654 142874 15706
rect 142874 15654 142876 15706
rect 142820 15652 142876 15654
rect 142924 15706 142980 15708
rect 142924 15654 142926 15706
rect 142926 15654 142978 15706
rect 142978 15654 142980 15706
rect 142924 15652 142980 15654
rect 142716 14138 142772 14140
rect 142716 14086 142718 14138
rect 142718 14086 142770 14138
rect 142770 14086 142772 14138
rect 142716 14084 142772 14086
rect 142820 14138 142876 14140
rect 142820 14086 142822 14138
rect 142822 14086 142874 14138
rect 142874 14086 142876 14138
rect 142820 14084 142876 14086
rect 142924 14138 142980 14140
rect 142924 14086 142926 14138
rect 142926 14086 142978 14138
rect 142978 14086 142980 14138
rect 142924 14084 142980 14086
rect 143612 12908 143668 12964
rect 142716 12570 142772 12572
rect 142716 12518 142718 12570
rect 142718 12518 142770 12570
rect 142770 12518 142772 12570
rect 142716 12516 142772 12518
rect 142820 12570 142876 12572
rect 142820 12518 142822 12570
rect 142822 12518 142874 12570
rect 142874 12518 142876 12570
rect 142820 12516 142876 12518
rect 142924 12570 142980 12572
rect 142924 12518 142926 12570
rect 142926 12518 142978 12570
rect 142978 12518 142980 12570
rect 142924 12516 142980 12518
rect 142716 11002 142772 11004
rect 142716 10950 142718 11002
rect 142718 10950 142770 11002
rect 142770 10950 142772 11002
rect 142716 10948 142772 10950
rect 142820 11002 142876 11004
rect 142820 10950 142822 11002
rect 142822 10950 142874 11002
rect 142874 10950 142876 11002
rect 142820 10948 142876 10950
rect 142924 11002 142980 11004
rect 142924 10950 142926 11002
rect 142926 10950 142978 11002
rect 142978 10950 142980 11002
rect 142924 10948 142980 10950
rect 142716 9434 142772 9436
rect 142716 9382 142718 9434
rect 142718 9382 142770 9434
rect 142770 9382 142772 9434
rect 142716 9380 142772 9382
rect 142820 9434 142876 9436
rect 142820 9382 142822 9434
rect 142822 9382 142874 9434
rect 142874 9382 142876 9434
rect 142820 9380 142876 9382
rect 142924 9434 142980 9436
rect 142924 9382 142926 9434
rect 142926 9382 142978 9434
rect 142978 9382 142980 9434
rect 142924 9380 142980 9382
rect 141932 9212 141988 9268
rect 142156 8146 142212 8148
rect 142156 8094 142158 8146
rect 142158 8094 142210 8146
rect 142210 8094 142212 8146
rect 142156 8092 142212 8094
rect 142716 7866 142772 7868
rect 142716 7814 142718 7866
rect 142718 7814 142770 7866
rect 142770 7814 142772 7866
rect 142716 7812 142772 7814
rect 142820 7866 142876 7868
rect 142820 7814 142822 7866
rect 142822 7814 142874 7866
rect 142874 7814 142876 7866
rect 142820 7812 142876 7814
rect 142924 7866 142980 7868
rect 142924 7814 142926 7866
rect 142926 7814 142978 7866
rect 142978 7814 142980 7866
rect 142924 7812 142980 7814
rect 142940 7644 142996 7700
rect 143276 7644 143332 7700
rect 141820 6412 141876 6468
rect 141820 5628 141876 5684
rect 141820 5404 141876 5460
rect 142492 6690 142548 6692
rect 142492 6638 142494 6690
rect 142494 6638 142546 6690
rect 142546 6638 142548 6690
rect 142492 6636 142548 6638
rect 142716 6298 142772 6300
rect 142716 6246 142718 6298
rect 142718 6246 142770 6298
rect 142770 6246 142772 6298
rect 142716 6244 142772 6246
rect 142820 6298 142876 6300
rect 142820 6246 142822 6298
rect 142822 6246 142874 6298
rect 142874 6246 142876 6298
rect 142820 6244 142876 6246
rect 142924 6298 142980 6300
rect 142924 6246 142926 6298
rect 142926 6246 142978 6298
rect 142978 6246 142980 6298
rect 142924 6244 142980 6246
rect 141932 5292 141988 5348
rect 142492 5180 142548 5236
rect 142268 5068 142324 5124
rect 141484 4956 141540 5012
rect 141260 4284 141316 4340
rect 143052 5122 143108 5124
rect 143052 5070 143054 5122
rect 143054 5070 143106 5122
rect 143106 5070 143108 5122
rect 143052 5068 143108 5070
rect 142716 4730 142772 4732
rect 142716 4678 142718 4730
rect 142718 4678 142770 4730
rect 142770 4678 142772 4730
rect 142716 4676 142772 4678
rect 142820 4730 142876 4732
rect 142820 4678 142822 4730
rect 142822 4678 142874 4730
rect 142874 4678 142876 4730
rect 142820 4676 142876 4678
rect 142924 4730 142980 4732
rect 142924 4678 142926 4730
rect 142926 4678 142978 4730
rect 142978 4678 142980 4730
rect 142924 4676 142980 4678
rect 143500 4338 143556 4340
rect 143500 4286 143502 4338
rect 143502 4286 143554 4338
rect 143554 4286 143556 4338
rect 143500 4284 143556 4286
rect 143052 4226 143108 4228
rect 143052 4174 143054 4226
rect 143054 4174 143106 4226
rect 143106 4174 143108 4226
rect 143052 4172 143108 4174
rect 142828 3666 142884 3668
rect 142828 3614 142830 3666
rect 142830 3614 142882 3666
rect 142882 3614 142884 3666
rect 142828 3612 142884 3614
rect 144060 7474 144116 7476
rect 144060 7422 144062 7474
rect 144062 7422 144114 7474
rect 144114 7422 144116 7474
rect 144060 7420 144116 7422
rect 145180 7084 145236 7140
rect 145292 7980 145348 8036
rect 145180 6860 145236 6916
rect 145068 6748 145124 6804
rect 144620 6578 144676 6580
rect 144620 6526 144622 6578
rect 144622 6526 144674 6578
rect 144674 6526 144676 6578
rect 144620 6524 144676 6526
rect 144284 6466 144340 6468
rect 144284 6414 144286 6466
rect 144286 6414 144338 6466
rect 144338 6414 144340 6466
rect 144284 6412 144340 6414
rect 143612 3612 143668 3668
rect 142716 3162 142772 3164
rect 142716 3110 142718 3162
rect 142718 3110 142770 3162
rect 142770 3110 142772 3162
rect 142716 3108 142772 3110
rect 142820 3162 142876 3164
rect 142820 3110 142822 3162
rect 142822 3110 142874 3162
rect 142874 3110 142876 3162
rect 142820 3108 142876 3110
rect 142924 3162 142980 3164
rect 142924 3110 142926 3162
rect 142926 3110 142978 3162
rect 142978 3110 142980 3162
rect 142924 3108 142980 3110
rect 141036 2604 141092 2660
rect 144284 5628 144340 5684
rect 144956 5122 145012 5124
rect 144956 5070 144958 5122
rect 144958 5070 145010 5122
rect 145010 5070 145012 5122
rect 144956 5068 145012 5070
rect 145740 7644 145796 7700
rect 145404 7084 145460 7140
rect 148204 13468 148260 13524
rect 146412 12796 146468 12852
rect 146188 10444 146244 10500
rect 146076 9436 146132 9492
rect 145852 6690 145908 6692
rect 145852 6638 145854 6690
rect 145854 6638 145906 6690
rect 145906 6638 145908 6690
rect 145852 6636 145908 6638
rect 147756 11676 147812 11732
rect 146860 11506 146916 11508
rect 146860 11454 146862 11506
rect 146862 11454 146914 11506
rect 146914 11454 146916 11506
rect 146860 11452 146916 11454
rect 147308 11506 147364 11508
rect 147308 11454 147310 11506
rect 147310 11454 147362 11506
rect 147362 11454 147364 11506
rect 147308 11452 147364 11454
rect 147532 10498 147588 10500
rect 147532 10446 147534 10498
rect 147534 10446 147586 10498
rect 147586 10446 147588 10498
rect 147532 10444 147588 10446
rect 145740 5516 145796 5572
rect 145404 5404 145460 5460
rect 144508 4172 144564 4228
rect 147644 6972 147700 7028
rect 158076 46282 158132 46284
rect 158076 46230 158078 46282
rect 158078 46230 158130 46282
rect 158130 46230 158132 46282
rect 158076 46228 158132 46230
rect 158180 46282 158236 46284
rect 158180 46230 158182 46282
rect 158182 46230 158234 46282
rect 158234 46230 158236 46282
rect 158180 46228 158236 46230
rect 158284 46282 158340 46284
rect 158284 46230 158286 46282
rect 158286 46230 158338 46282
rect 158338 46230 158340 46282
rect 158284 46228 158340 46230
rect 172508 45836 172564 45892
rect 173292 45890 173348 45892
rect 173292 45838 173294 45890
rect 173294 45838 173346 45890
rect 173346 45838 173348 45890
rect 173292 45836 173348 45838
rect 176316 45836 176372 45892
rect 177100 45890 177156 45892
rect 177100 45838 177102 45890
rect 177102 45838 177154 45890
rect 177154 45838 177156 45890
rect 177100 45836 177156 45838
rect 188796 46282 188852 46284
rect 188796 46230 188798 46282
rect 188798 46230 188850 46282
rect 188850 46230 188852 46282
rect 188796 46228 188852 46230
rect 188900 46282 188956 46284
rect 188900 46230 188902 46282
rect 188902 46230 188954 46282
rect 188954 46230 188956 46282
rect 188900 46228 188956 46230
rect 189004 46282 189060 46284
rect 189004 46230 189006 46282
rect 189006 46230 189058 46282
rect 189058 46230 189060 46282
rect 189004 46228 189060 46230
rect 184044 45836 184100 45892
rect 184828 45890 184884 45892
rect 184828 45838 184830 45890
rect 184830 45838 184882 45890
rect 184882 45838 184884 45890
rect 184828 45836 184884 45838
rect 187292 45724 187348 45780
rect 152124 45276 152180 45332
rect 152124 44994 152180 44996
rect 152124 44942 152126 44994
rect 152126 44942 152178 44994
rect 152178 44942 152180 44994
rect 152124 44940 152180 44942
rect 153356 45330 153412 45332
rect 153356 45278 153358 45330
rect 153358 45278 153410 45330
rect 153410 45278 153412 45330
rect 153356 45276 153412 45278
rect 158076 44714 158132 44716
rect 158076 44662 158078 44714
rect 158078 44662 158130 44714
rect 158130 44662 158132 44714
rect 158076 44660 158132 44662
rect 158180 44714 158236 44716
rect 158180 44662 158182 44714
rect 158182 44662 158234 44714
rect 158234 44662 158236 44714
rect 158180 44660 158236 44662
rect 158284 44714 158340 44716
rect 158284 44662 158286 44714
rect 158286 44662 158338 44714
rect 158338 44662 158340 44714
rect 158284 44660 158340 44662
rect 153244 12684 153300 12740
rect 153692 14252 153748 14308
rect 150332 11676 150388 11732
rect 150780 12572 150836 12628
rect 149212 11506 149268 11508
rect 149212 11454 149214 11506
rect 149214 11454 149266 11506
rect 149266 11454 149268 11506
rect 149212 11452 149268 11454
rect 147868 10834 147924 10836
rect 147868 10782 147870 10834
rect 147870 10782 147922 10834
rect 147922 10782 147924 10834
rect 147868 10780 147924 10782
rect 148204 10780 148260 10836
rect 148204 10444 148260 10500
rect 148764 9772 148820 9828
rect 150668 11452 150724 11508
rect 149660 10610 149716 10612
rect 149660 10558 149662 10610
rect 149662 10558 149714 10610
rect 149714 10558 149716 10610
rect 149660 10556 149716 10558
rect 148876 10220 148932 10276
rect 147868 8370 147924 8372
rect 147868 8318 147870 8370
rect 147870 8318 147922 8370
rect 147922 8318 147924 8370
rect 147868 8316 147924 8318
rect 147980 9548 148036 9604
rect 147868 7698 147924 7700
rect 147868 7646 147870 7698
rect 147870 7646 147922 7698
rect 147922 7646 147924 7698
rect 147868 7644 147924 7646
rect 148652 9602 148708 9604
rect 148652 9550 148654 9602
rect 148654 9550 148706 9602
rect 148706 9550 148708 9602
rect 148652 9548 148708 9550
rect 148428 9266 148484 9268
rect 148428 9214 148430 9266
rect 148430 9214 148482 9266
rect 148482 9214 148484 9266
rect 148428 9212 148484 9214
rect 148540 9154 148596 9156
rect 148540 9102 148542 9154
rect 148542 9102 148594 9154
rect 148594 9102 148596 9154
rect 148540 9100 148596 9102
rect 148540 8370 148596 8372
rect 148540 8318 148542 8370
rect 148542 8318 148594 8370
rect 148594 8318 148596 8370
rect 148540 8316 148596 8318
rect 149324 9100 149380 9156
rect 149548 9772 149604 9828
rect 150108 9772 150164 9828
rect 149772 9212 149828 9268
rect 149660 8930 149716 8932
rect 149660 8878 149662 8930
rect 149662 8878 149714 8930
rect 149714 8878 149716 8930
rect 149660 8876 149716 8878
rect 146076 5740 146132 5796
rect 145852 5234 145908 5236
rect 145852 5182 145854 5234
rect 145854 5182 145906 5234
rect 145906 5182 145908 5234
rect 145852 5180 145908 5182
rect 148092 6748 148148 6804
rect 147308 5852 147364 5908
rect 146636 5068 146692 5124
rect 146076 3612 146132 3668
rect 144508 2156 144564 2212
rect 144396 1596 144452 1652
rect 145404 1372 145460 1428
rect 146860 4898 146916 4900
rect 146860 4846 146862 4898
rect 146862 4846 146914 4898
rect 146914 4846 146916 4898
rect 146860 4844 146916 4846
rect 147084 4338 147140 4340
rect 147084 4286 147086 4338
rect 147086 4286 147138 4338
rect 147138 4286 147140 4338
rect 147084 4284 147140 4286
rect 147420 4956 147476 5012
rect 150108 9436 150164 9492
rect 150556 10220 150612 10276
rect 150668 9548 150724 9604
rect 151228 10610 151284 10612
rect 151228 10558 151230 10610
rect 151230 10558 151282 10610
rect 151282 10558 151284 10610
rect 151228 10556 151284 10558
rect 150780 9436 150836 9492
rect 151452 10108 151508 10164
rect 151116 9212 151172 9268
rect 151564 9826 151620 9828
rect 151564 9774 151566 9826
rect 151566 9774 151618 9826
rect 151618 9774 151620 9826
rect 151564 9772 151620 9774
rect 151676 9548 151732 9604
rect 151004 8204 151060 8260
rect 148204 7420 148260 7476
rect 148764 7420 148820 7476
rect 148876 7308 148932 7364
rect 148540 5516 148596 5572
rect 147420 4172 147476 4228
rect 148316 4284 148372 4340
rect 148540 5068 148596 5124
rect 148988 6412 149044 6468
rect 149100 5794 149156 5796
rect 149100 5742 149102 5794
rect 149102 5742 149154 5794
rect 149154 5742 149156 5794
rect 149100 5740 149156 5742
rect 149100 4562 149156 4564
rect 149100 4510 149102 4562
rect 149102 4510 149154 4562
rect 149154 4510 149156 4562
rect 149100 4508 149156 4510
rect 147308 2380 147364 2436
rect 148652 3612 148708 3668
rect 148316 2380 148372 2436
rect 149996 7196 150052 7252
rect 150220 7084 150276 7140
rect 150108 6972 150164 7028
rect 152124 9212 152180 9268
rect 152236 10332 152292 10388
rect 151676 8428 151732 8484
rect 149660 6188 149716 6244
rect 149436 5906 149492 5908
rect 149436 5854 149438 5906
rect 149438 5854 149490 5906
rect 149490 5854 149492 5906
rect 149436 5852 149492 5854
rect 149884 6018 149940 6020
rect 149884 5966 149886 6018
rect 149886 5966 149938 6018
rect 149938 5966 149940 6018
rect 149884 5964 149940 5966
rect 150108 5906 150164 5908
rect 150108 5854 150110 5906
rect 150110 5854 150162 5906
rect 150162 5854 150164 5906
rect 150108 5852 150164 5854
rect 149772 4508 149828 4564
rect 150220 5794 150276 5796
rect 150220 5742 150222 5794
rect 150222 5742 150274 5794
rect 150274 5742 150276 5794
rect 150220 5740 150276 5742
rect 150332 5628 150388 5684
rect 150668 5852 150724 5908
rect 150556 5516 150612 5572
rect 150332 4844 150388 4900
rect 150892 7474 150948 7476
rect 150892 7422 150894 7474
rect 150894 7422 150946 7474
rect 150946 7422 150948 7474
rect 150892 7420 150948 7422
rect 150780 4732 150836 4788
rect 151116 7308 151172 7364
rect 151228 7420 151284 7476
rect 151116 6690 151172 6692
rect 151116 6638 151118 6690
rect 151118 6638 151170 6690
rect 151170 6638 151172 6690
rect 151116 6636 151172 6638
rect 151452 6860 151508 6916
rect 151452 6188 151508 6244
rect 153132 10220 153188 10276
rect 153580 10498 153636 10500
rect 153580 10446 153582 10498
rect 153582 10446 153634 10498
rect 153634 10446 153636 10498
rect 153580 10444 153636 10446
rect 153244 9884 153300 9940
rect 152460 8988 152516 9044
rect 152348 8258 152404 8260
rect 152348 8206 152350 8258
rect 152350 8206 152402 8258
rect 152402 8206 152404 8258
rect 152348 8204 152404 8206
rect 152796 8428 152852 8484
rect 151900 7756 151956 7812
rect 152124 7474 152180 7476
rect 152124 7422 152126 7474
rect 152126 7422 152178 7474
rect 152178 7422 152180 7474
rect 152124 7420 152180 7422
rect 152236 7308 152292 7364
rect 152124 7084 152180 7140
rect 151340 5906 151396 5908
rect 151340 5854 151342 5906
rect 151342 5854 151394 5906
rect 151394 5854 151396 5906
rect 151340 5852 151396 5854
rect 151228 4956 151284 5012
rect 152124 5964 152180 6020
rect 151900 5852 151956 5908
rect 150220 4450 150276 4452
rect 150220 4398 150222 4450
rect 150222 4398 150274 4450
rect 150274 4398 150276 4450
rect 150220 4396 150276 4398
rect 149436 3948 149492 4004
rect 150332 3948 150388 4004
rect 151452 3836 151508 3892
rect 152012 3724 152068 3780
rect 151340 3388 151396 3444
rect 151452 3500 151508 3556
rect 151228 2268 151284 2324
rect 149212 1484 149268 1540
rect 152908 7474 152964 7476
rect 152908 7422 152910 7474
rect 152910 7422 152962 7474
rect 152962 7422 152964 7474
rect 152908 7420 152964 7422
rect 152460 7362 152516 7364
rect 152460 7310 152462 7362
rect 152462 7310 152514 7362
rect 152514 7310 152516 7362
rect 152460 7308 152516 7310
rect 152684 6300 152740 6356
rect 152572 6188 152628 6244
rect 152460 6076 152516 6132
rect 153244 8428 153300 8484
rect 153132 7756 153188 7812
rect 153468 8764 153524 8820
rect 153244 6412 153300 6468
rect 152796 5180 152852 5236
rect 152460 5010 152516 5012
rect 152460 4958 152462 5010
rect 152462 4958 152514 5010
rect 152514 4958 152516 5010
rect 152460 4956 152516 4958
rect 152572 4620 152628 4676
rect 152460 3836 152516 3892
rect 152796 3666 152852 3668
rect 152796 3614 152798 3666
rect 152798 3614 152850 3666
rect 152850 3614 152852 3666
rect 152796 3612 152852 3614
rect 152572 3388 152628 3444
rect 153020 5346 153076 5348
rect 153020 5294 153022 5346
rect 153022 5294 153074 5346
rect 153074 5294 153076 5346
rect 153020 5292 153076 5294
rect 153244 4844 153300 4900
rect 154588 12684 154644 12740
rect 154028 10668 154084 10724
rect 155148 10892 155204 10948
rect 154924 10722 154980 10724
rect 154924 10670 154926 10722
rect 154926 10670 154978 10722
rect 154978 10670 154980 10722
rect 154924 10668 154980 10670
rect 154812 10220 154868 10276
rect 155596 10444 155652 10500
rect 155596 9996 155652 10052
rect 153916 9042 153972 9044
rect 153916 8990 153918 9042
rect 153918 8990 153970 9042
rect 153970 8990 153972 9042
rect 153916 8988 153972 8990
rect 153804 8428 153860 8484
rect 153580 7420 153636 7476
rect 156492 11452 156548 11508
rect 156044 11340 156100 11396
rect 156044 9772 156100 9828
rect 156268 9772 156324 9828
rect 155708 9602 155764 9604
rect 155708 9550 155710 9602
rect 155710 9550 155762 9602
rect 155762 9550 155764 9602
rect 155708 9548 155764 9550
rect 155372 8428 155428 8484
rect 155148 7644 155204 7700
rect 154252 6860 154308 6916
rect 153692 5852 153748 5908
rect 153692 4172 153748 4228
rect 153580 3836 153636 3892
rect 153356 3554 153412 3556
rect 153356 3502 153358 3554
rect 153358 3502 153410 3554
rect 153410 3502 153412 3554
rect 153356 3500 153412 3502
rect 154028 6076 154084 6132
rect 153916 5404 153972 5460
rect 154924 7308 154980 7364
rect 154700 6636 154756 6692
rect 153916 5180 153972 5236
rect 153916 4508 153972 4564
rect 154812 5964 154868 6020
rect 154700 5068 154756 5124
rect 154924 5404 154980 5460
rect 154812 4898 154868 4900
rect 154812 4846 154814 4898
rect 154814 4846 154866 4898
rect 154866 4846 154868 4898
rect 154812 4844 154868 4846
rect 155148 7196 155204 7252
rect 156044 9266 156100 9268
rect 156044 9214 156046 9266
rect 156046 9214 156098 9266
rect 156098 9214 156100 9266
rect 156044 9212 156100 9214
rect 155820 6860 155876 6916
rect 156044 6412 156100 6468
rect 155932 5404 155988 5460
rect 155820 5292 155876 5348
rect 155820 5068 155876 5124
rect 155036 4620 155092 4676
rect 155260 4562 155316 4564
rect 155260 4510 155262 4562
rect 155262 4510 155314 4562
rect 155314 4510 155316 4562
rect 155260 4508 155316 4510
rect 154140 4172 154196 4228
rect 154476 3836 154532 3892
rect 154140 3388 154196 3444
rect 152908 2492 152964 2548
rect 155036 3388 155092 3444
rect 155708 3554 155764 3556
rect 155708 3502 155710 3554
rect 155710 3502 155762 3554
rect 155762 3502 155764 3554
rect 155708 3500 155764 3502
rect 157164 11564 157220 11620
rect 156716 11394 156772 11396
rect 156716 11342 156718 11394
rect 156718 11342 156770 11394
rect 156770 11342 156772 11394
rect 156716 11340 156772 11342
rect 156716 11004 156772 11060
rect 156940 10892 156996 10948
rect 156716 10444 156772 10500
rect 157164 9996 157220 10052
rect 156828 9826 156884 9828
rect 156828 9774 156830 9826
rect 156830 9774 156882 9826
rect 156882 9774 156884 9826
rect 156828 9772 156884 9774
rect 157052 9714 157108 9716
rect 157052 9662 157054 9714
rect 157054 9662 157106 9714
rect 157106 9662 157108 9714
rect 157052 9660 157108 9662
rect 156380 8092 156436 8148
rect 156604 7196 156660 7252
rect 158076 43146 158132 43148
rect 158076 43094 158078 43146
rect 158078 43094 158130 43146
rect 158130 43094 158132 43146
rect 158076 43092 158132 43094
rect 158180 43146 158236 43148
rect 158180 43094 158182 43146
rect 158182 43094 158234 43146
rect 158234 43094 158236 43146
rect 158180 43092 158236 43094
rect 158284 43146 158340 43148
rect 158284 43094 158286 43146
rect 158286 43094 158338 43146
rect 158338 43094 158340 43146
rect 158284 43092 158340 43094
rect 158076 41578 158132 41580
rect 158076 41526 158078 41578
rect 158078 41526 158130 41578
rect 158130 41526 158132 41578
rect 158076 41524 158132 41526
rect 158180 41578 158236 41580
rect 158180 41526 158182 41578
rect 158182 41526 158234 41578
rect 158234 41526 158236 41578
rect 158180 41524 158236 41526
rect 158284 41578 158340 41580
rect 158284 41526 158286 41578
rect 158286 41526 158338 41578
rect 158338 41526 158340 41578
rect 158284 41524 158340 41526
rect 158076 40010 158132 40012
rect 158076 39958 158078 40010
rect 158078 39958 158130 40010
rect 158130 39958 158132 40010
rect 158076 39956 158132 39958
rect 158180 40010 158236 40012
rect 158180 39958 158182 40010
rect 158182 39958 158234 40010
rect 158234 39958 158236 40010
rect 158180 39956 158236 39958
rect 158284 40010 158340 40012
rect 158284 39958 158286 40010
rect 158286 39958 158338 40010
rect 158338 39958 158340 40010
rect 158284 39956 158340 39958
rect 158076 38442 158132 38444
rect 158076 38390 158078 38442
rect 158078 38390 158130 38442
rect 158130 38390 158132 38442
rect 158076 38388 158132 38390
rect 158180 38442 158236 38444
rect 158180 38390 158182 38442
rect 158182 38390 158234 38442
rect 158234 38390 158236 38442
rect 158180 38388 158236 38390
rect 158284 38442 158340 38444
rect 158284 38390 158286 38442
rect 158286 38390 158338 38442
rect 158338 38390 158340 38442
rect 158284 38388 158340 38390
rect 158076 36874 158132 36876
rect 158076 36822 158078 36874
rect 158078 36822 158130 36874
rect 158130 36822 158132 36874
rect 158076 36820 158132 36822
rect 158180 36874 158236 36876
rect 158180 36822 158182 36874
rect 158182 36822 158234 36874
rect 158234 36822 158236 36874
rect 158180 36820 158236 36822
rect 158284 36874 158340 36876
rect 158284 36822 158286 36874
rect 158286 36822 158338 36874
rect 158338 36822 158340 36874
rect 158284 36820 158340 36822
rect 158076 35306 158132 35308
rect 158076 35254 158078 35306
rect 158078 35254 158130 35306
rect 158130 35254 158132 35306
rect 158076 35252 158132 35254
rect 158180 35306 158236 35308
rect 158180 35254 158182 35306
rect 158182 35254 158234 35306
rect 158234 35254 158236 35306
rect 158180 35252 158236 35254
rect 158284 35306 158340 35308
rect 158284 35254 158286 35306
rect 158286 35254 158338 35306
rect 158338 35254 158340 35306
rect 158284 35252 158340 35254
rect 158076 33738 158132 33740
rect 158076 33686 158078 33738
rect 158078 33686 158130 33738
rect 158130 33686 158132 33738
rect 158076 33684 158132 33686
rect 158180 33738 158236 33740
rect 158180 33686 158182 33738
rect 158182 33686 158234 33738
rect 158234 33686 158236 33738
rect 158180 33684 158236 33686
rect 158284 33738 158340 33740
rect 158284 33686 158286 33738
rect 158286 33686 158338 33738
rect 158338 33686 158340 33738
rect 158284 33684 158340 33686
rect 158076 32170 158132 32172
rect 158076 32118 158078 32170
rect 158078 32118 158130 32170
rect 158130 32118 158132 32170
rect 158076 32116 158132 32118
rect 158180 32170 158236 32172
rect 158180 32118 158182 32170
rect 158182 32118 158234 32170
rect 158234 32118 158236 32170
rect 158180 32116 158236 32118
rect 158284 32170 158340 32172
rect 158284 32118 158286 32170
rect 158286 32118 158338 32170
rect 158338 32118 158340 32170
rect 158284 32116 158340 32118
rect 158076 30602 158132 30604
rect 158076 30550 158078 30602
rect 158078 30550 158130 30602
rect 158130 30550 158132 30602
rect 158076 30548 158132 30550
rect 158180 30602 158236 30604
rect 158180 30550 158182 30602
rect 158182 30550 158234 30602
rect 158234 30550 158236 30602
rect 158180 30548 158236 30550
rect 158284 30602 158340 30604
rect 158284 30550 158286 30602
rect 158286 30550 158338 30602
rect 158338 30550 158340 30602
rect 158284 30548 158340 30550
rect 158076 29034 158132 29036
rect 158076 28982 158078 29034
rect 158078 28982 158130 29034
rect 158130 28982 158132 29034
rect 158076 28980 158132 28982
rect 158180 29034 158236 29036
rect 158180 28982 158182 29034
rect 158182 28982 158234 29034
rect 158234 28982 158236 29034
rect 158180 28980 158236 28982
rect 158284 29034 158340 29036
rect 158284 28982 158286 29034
rect 158286 28982 158338 29034
rect 158338 28982 158340 29034
rect 158284 28980 158340 28982
rect 158076 27466 158132 27468
rect 158076 27414 158078 27466
rect 158078 27414 158130 27466
rect 158130 27414 158132 27466
rect 158076 27412 158132 27414
rect 158180 27466 158236 27468
rect 158180 27414 158182 27466
rect 158182 27414 158234 27466
rect 158234 27414 158236 27466
rect 158180 27412 158236 27414
rect 158284 27466 158340 27468
rect 158284 27414 158286 27466
rect 158286 27414 158338 27466
rect 158338 27414 158340 27466
rect 158284 27412 158340 27414
rect 158076 25898 158132 25900
rect 158076 25846 158078 25898
rect 158078 25846 158130 25898
rect 158130 25846 158132 25898
rect 158076 25844 158132 25846
rect 158180 25898 158236 25900
rect 158180 25846 158182 25898
rect 158182 25846 158234 25898
rect 158234 25846 158236 25898
rect 158180 25844 158236 25846
rect 158284 25898 158340 25900
rect 158284 25846 158286 25898
rect 158286 25846 158338 25898
rect 158338 25846 158340 25898
rect 158284 25844 158340 25846
rect 158076 24330 158132 24332
rect 158076 24278 158078 24330
rect 158078 24278 158130 24330
rect 158130 24278 158132 24330
rect 158076 24276 158132 24278
rect 158180 24330 158236 24332
rect 158180 24278 158182 24330
rect 158182 24278 158234 24330
rect 158234 24278 158236 24330
rect 158180 24276 158236 24278
rect 158284 24330 158340 24332
rect 158284 24278 158286 24330
rect 158286 24278 158338 24330
rect 158338 24278 158340 24330
rect 158284 24276 158340 24278
rect 158076 22762 158132 22764
rect 158076 22710 158078 22762
rect 158078 22710 158130 22762
rect 158130 22710 158132 22762
rect 158076 22708 158132 22710
rect 158180 22762 158236 22764
rect 158180 22710 158182 22762
rect 158182 22710 158234 22762
rect 158234 22710 158236 22762
rect 158180 22708 158236 22710
rect 158284 22762 158340 22764
rect 158284 22710 158286 22762
rect 158286 22710 158338 22762
rect 158338 22710 158340 22762
rect 158284 22708 158340 22710
rect 158076 21194 158132 21196
rect 158076 21142 158078 21194
rect 158078 21142 158130 21194
rect 158130 21142 158132 21194
rect 158076 21140 158132 21142
rect 158180 21194 158236 21196
rect 158180 21142 158182 21194
rect 158182 21142 158234 21194
rect 158234 21142 158236 21194
rect 158180 21140 158236 21142
rect 158284 21194 158340 21196
rect 158284 21142 158286 21194
rect 158286 21142 158338 21194
rect 158338 21142 158340 21194
rect 158284 21140 158340 21142
rect 158076 19626 158132 19628
rect 158076 19574 158078 19626
rect 158078 19574 158130 19626
rect 158130 19574 158132 19626
rect 158076 19572 158132 19574
rect 158180 19626 158236 19628
rect 158180 19574 158182 19626
rect 158182 19574 158234 19626
rect 158234 19574 158236 19626
rect 158180 19572 158236 19574
rect 158284 19626 158340 19628
rect 158284 19574 158286 19626
rect 158286 19574 158338 19626
rect 158338 19574 158340 19626
rect 158284 19572 158340 19574
rect 158076 18058 158132 18060
rect 158076 18006 158078 18058
rect 158078 18006 158130 18058
rect 158130 18006 158132 18058
rect 158076 18004 158132 18006
rect 158180 18058 158236 18060
rect 158180 18006 158182 18058
rect 158182 18006 158234 18058
rect 158234 18006 158236 18058
rect 158180 18004 158236 18006
rect 158284 18058 158340 18060
rect 158284 18006 158286 18058
rect 158286 18006 158338 18058
rect 158338 18006 158340 18058
rect 158284 18004 158340 18006
rect 158076 16490 158132 16492
rect 158076 16438 158078 16490
rect 158078 16438 158130 16490
rect 158130 16438 158132 16490
rect 158076 16436 158132 16438
rect 158180 16490 158236 16492
rect 158180 16438 158182 16490
rect 158182 16438 158234 16490
rect 158234 16438 158236 16490
rect 158180 16436 158236 16438
rect 158284 16490 158340 16492
rect 158284 16438 158286 16490
rect 158286 16438 158338 16490
rect 158338 16438 158340 16490
rect 158284 16436 158340 16438
rect 158076 14922 158132 14924
rect 158076 14870 158078 14922
rect 158078 14870 158130 14922
rect 158130 14870 158132 14922
rect 158076 14868 158132 14870
rect 158180 14922 158236 14924
rect 158180 14870 158182 14922
rect 158182 14870 158234 14922
rect 158234 14870 158236 14922
rect 158180 14868 158236 14870
rect 158284 14922 158340 14924
rect 158284 14870 158286 14922
rect 158286 14870 158338 14922
rect 158338 14870 158340 14922
rect 158284 14868 158340 14870
rect 158076 13354 158132 13356
rect 158076 13302 158078 13354
rect 158078 13302 158130 13354
rect 158130 13302 158132 13354
rect 158076 13300 158132 13302
rect 158180 13354 158236 13356
rect 158180 13302 158182 13354
rect 158182 13302 158234 13354
rect 158234 13302 158236 13354
rect 158180 13300 158236 13302
rect 158284 13354 158340 13356
rect 158284 13302 158286 13354
rect 158286 13302 158338 13354
rect 158338 13302 158340 13354
rect 158284 13300 158340 13302
rect 158076 11786 158132 11788
rect 158076 11734 158078 11786
rect 158078 11734 158130 11786
rect 158130 11734 158132 11786
rect 158076 11732 158132 11734
rect 158180 11786 158236 11788
rect 158180 11734 158182 11786
rect 158182 11734 158234 11786
rect 158234 11734 158236 11786
rect 158180 11732 158236 11734
rect 158284 11786 158340 11788
rect 158284 11734 158286 11786
rect 158286 11734 158338 11786
rect 158338 11734 158340 11786
rect 158284 11732 158340 11734
rect 157724 11564 157780 11620
rect 160300 11452 160356 11508
rect 159852 11116 159908 11172
rect 158076 10218 158132 10220
rect 158076 10166 158078 10218
rect 158078 10166 158130 10218
rect 158130 10166 158132 10218
rect 158076 10164 158132 10166
rect 158180 10218 158236 10220
rect 158180 10166 158182 10218
rect 158182 10166 158234 10218
rect 158234 10166 158236 10218
rect 158180 10164 158236 10166
rect 158284 10218 158340 10220
rect 158284 10166 158286 10218
rect 158286 10166 158338 10218
rect 158338 10166 158340 10218
rect 158284 10164 158340 10166
rect 157276 9602 157332 9604
rect 157276 9550 157278 9602
rect 157278 9550 157330 9602
rect 157330 9550 157332 9602
rect 157276 9548 157332 9550
rect 156828 8764 156884 8820
rect 158076 8650 158132 8652
rect 158076 8598 158078 8650
rect 158078 8598 158130 8650
rect 158130 8598 158132 8650
rect 158076 8596 158132 8598
rect 158180 8650 158236 8652
rect 158180 8598 158182 8650
rect 158182 8598 158234 8650
rect 158234 8598 158236 8650
rect 158180 8596 158236 8598
rect 158284 8650 158340 8652
rect 158284 8598 158286 8650
rect 158286 8598 158338 8650
rect 158338 8598 158340 8650
rect 158284 8596 158340 8598
rect 156828 8316 156884 8372
rect 159292 8204 159348 8260
rect 158076 7082 158132 7084
rect 158076 7030 158078 7082
rect 158078 7030 158130 7082
rect 158130 7030 158132 7082
rect 158076 7028 158132 7030
rect 158180 7082 158236 7084
rect 158180 7030 158182 7082
rect 158182 7030 158234 7082
rect 158234 7030 158236 7082
rect 158180 7028 158236 7030
rect 158284 7082 158340 7084
rect 158284 7030 158286 7082
rect 158286 7030 158338 7082
rect 158338 7030 158340 7082
rect 158284 7028 158340 7030
rect 156828 6130 156884 6132
rect 156828 6078 156830 6130
rect 156830 6078 156882 6130
rect 156882 6078 156884 6130
rect 156828 6076 156884 6078
rect 157948 6130 158004 6132
rect 157948 6078 157950 6130
rect 157950 6078 158002 6130
rect 158002 6078 158004 6130
rect 157948 6076 158004 6078
rect 159628 6636 159684 6692
rect 157724 5964 157780 6020
rect 157164 5628 157220 5684
rect 156828 5292 156884 5348
rect 156828 5068 156884 5124
rect 157388 5292 157444 5348
rect 157276 5180 157332 5236
rect 156268 4956 156324 5012
rect 156604 4956 156660 5012
rect 156044 3724 156100 3780
rect 155932 3500 155988 3556
rect 158076 5514 158132 5516
rect 158076 5462 158078 5514
rect 158078 5462 158130 5514
rect 158130 5462 158132 5514
rect 158076 5460 158132 5462
rect 158180 5514 158236 5516
rect 158180 5462 158182 5514
rect 158182 5462 158234 5514
rect 158234 5462 158236 5514
rect 158180 5460 158236 5462
rect 158284 5514 158340 5516
rect 158284 5462 158286 5514
rect 158286 5462 158338 5514
rect 158338 5462 158340 5514
rect 158284 5460 158340 5462
rect 157836 5292 157892 5348
rect 157948 5234 158004 5236
rect 157948 5182 157950 5234
rect 157950 5182 158002 5234
rect 158002 5182 158004 5234
rect 157948 5180 158004 5182
rect 159628 6412 159684 6468
rect 160300 10610 160356 10612
rect 160300 10558 160302 10610
rect 160302 10558 160354 10610
rect 160354 10558 160356 10610
rect 160300 10556 160356 10558
rect 160076 9436 160132 9492
rect 160076 7756 160132 7812
rect 160076 6524 160132 6580
rect 159964 6076 160020 6132
rect 162876 15932 162932 15988
rect 160748 11676 160804 11732
rect 160524 10722 160580 10724
rect 160524 10670 160526 10722
rect 160526 10670 160578 10722
rect 160578 10670 160580 10722
rect 160524 10668 160580 10670
rect 162876 11676 162932 11732
rect 163324 12066 163380 12068
rect 163324 12014 163326 12066
rect 163326 12014 163378 12066
rect 163378 12014 163380 12066
rect 163324 12012 163380 12014
rect 161980 10892 162036 10948
rect 161532 10834 161588 10836
rect 161532 10782 161534 10834
rect 161534 10782 161586 10834
rect 161586 10782 161588 10834
rect 161532 10780 161588 10782
rect 160412 10108 160468 10164
rect 161196 10610 161252 10612
rect 161196 10558 161198 10610
rect 161198 10558 161250 10610
rect 161250 10558 161252 10610
rect 161196 10556 161252 10558
rect 162092 10722 162148 10724
rect 162092 10670 162094 10722
rect 162094 10670 162146 10722
rect 162146 10670 162148 10722
rect 162092 10668 162148 10670
rect 161644 10444 161700 10500
rect 161532 9436 161588 9492
rect 160636 8876 160692 8932
rect 161196 8428 161252 8484
rect 160300 7308 160356 7364
rect 160300 6076 160356 6132
rect 160524 6748 160580 6804
rect 159740 5516 159796 5572
rect 159292 5068 159348 5124
rect 158284 5010 158340 5012
rect 158284 4958 158286 5010
rect 158286 4958 158338 5010
rect 158338 4958 158340 5010
rect 158284 4956 158340 4958
rect 161084 7362 161140 7364
rect 161084 7310 161086 7362
rect 161086 7310 161138 7362
rect 161138 7310 161140 7362
rect 161084 7308 161140 7310
rect 162652 11170 162708 11172
rect 162652 11118 162654 11170
rect 162654 11118 162706 11170
rect 162706 11118 162708 11170
rect 162652 11116 162708 11118
rect 162316 10834 162372 10836
rect 162316 10782 162318 10834
rect 162318 10782 162370 10834
rect 162370 10782 162372 10834
rect 162316 10780 162372 10782
rect 162540 10610 162596 10612
rect 162540 10558 162542 10610
rect 162542 10558 162594 10610
rect 162594 10558 162596 10610
rect 162540 10556 162596 10558
rect 161756 7586 161812 7588
rect 161756 7534 161758 7586
rect 161758 7534 161810 7586
rect 161810 7534 161812 7586
rect 161756 7532 161812 7534
rect 162204 7532 162260 7588
rect 161420 7308 161476 7364
rect 161644 7196 161700 7252
rect 160972 6690 161028 6692
rect 160972 6638 160974 6690
rect 160974 6638 161026 6690
rect 161026 6638 161028 6690
rect 160972 6636 161028 6638
rect 160748 6466 160804 6468
rect 160748 6414 160750 6466
rect 160750 6414 160802 6466
rect 160802 6414 160804 6466
rect 160748 6412 160804 6414
rect 160748 6076 160804 6132
rect 160748 5516 160804 5572
rect 160524 5122 160580 5124
rect 160524 5070 160526 5122
rect 160526 5070 160578 5122
rect 160578 5070 160580 5122
rect 160524 5068 160580 5070
rect 157724 4732 157780 4788
rect 157836 4844 157892 4900
rect 157388 3724 157444 3780
rect 156604 3442 156660 3444
rect 156604 3390 156606 3442
rect 156606 3390 156658 3442
rect 156658 3390 156660 3442
rect 156604 3388 156660 3390
rect 157388 3442 157444 3444
rect 157388 3390 157390 3442
rect 157390 3390 157442 3442
rect 157442 3390 157444 3442
rect 157388 3388 157444 3390
rect 156380 2604 156436 2660
rect 158060 4898 158116 4900
rect 158060 4846 158062 4898
rect 158062 4846 158114 4898
rect 158114 4846 158116 4898
rect 158060 4844 158116 4846
rect 159740 4844 159796 4900
rect 158076 3946 158132 3948
rect 158076 3894 158078 3946
rect 158078 3894 158130 3946
rect 158130 3894 158132 3946
rect 158076 3892 158132 3894
rect 158180 3946 158236 3948
rect 158180 3894 158182 3946
rect 158182 3894 158234 3946
rect 158234 3894 158236 3946
rect 158180 3892 158236 3894
rect 158284 3946 158340 3948
rect 158284 3894 158286 3946
rect 158286 3894 158338 3946
rect 158338 3894 158340 3946
rect 158284 3892 158340 3894
rect 158172 3442 158228 3444
rect 158172 3390 158174 3442
rect 158174 3390 158226 3442
rect 158226 3390 158228 3442
rect 158172 3388 158228 3390
rect 159516 3442 159572 3444
rect 159516 3390 159518 3442
rect 159518 3390 159570 3442
rect 159570 3390 159572 3442
rect 159516 3388 159572 3390
rect 161532 6802 161588 6804
rect 161532 6750 161534 6802
rect 161534 6750 161586 6802
rect 161586 6750 161588 6802
rect 161532 6748 161588 6750
rect 161196 6636 161252 6692
rect 161420 6578 161476 6580
rect 161420 6526 161422 6578
rect 161422 6526 161474 6578
rect 161474 6526 161476 6578
rect 161420 6524 161476 6526
rect 161644 6466 161700 6468
rect 161644 6414 161646 6466
rect 161646 6414 161698 6466
rect 161698 6414 161700 6466
rect 161644 6412 161700 6414
rect 160636 3724 160692 3780
rect 160076 3442 160132 3444
rect 160076 3390 160078 3442
rect 160078 3390 160130 3442
rect 160130 3390 160132 3442
rect 160076 3388 160132 3390
rect 161980 6300 162036 6356
rect 161756 5404 161812 5460
rect 161868 5740 161924 5796
rect 161980 5180 162036 5236
rect 161532 5122 161588 5124
rect 161532 5070 161534 5122
rect 161534 5070 161586 5122
rect 161586 5070 161588 5122
rect 161532 5068 161588 5070
rect 161420 4844 161476 4900
rect 161756 4508 161812 4564
rect 162428 8258 162484 8260
rect 162428 8206 162430 8258
rect 162430 8206 162482 8258
rect 162482 8206 162484 8258
rect 162428 8204 162484 8206
rect 162540 7474 162596 7476
rect 162540 7422 162542 7474
rect 162542 7422 162594 7474
rect 162594 7422 162596 7474
rect 162540 7420 162596 7422
rect 162988 11564 163044 11620
rect 162876 11004 162932 11060
rect 167132 43708 167188 43764
rect 164444 11788 164500 11844
rect 164668 14140 164724 14196
rect 163996 11394 164052 11396
rect 163996 11342 163998 11394
rect 163998 11342 164050 11394
rect 164050 11342 164052 11394
rect 163996 11340 164052 11342
rect 164668 11340 164724 11396
rect 162988 10892 163044 10948
rect 162764 8540 162820 8596
rect 162764 8034 162820 8036
rect 162764 7982 162766 8034
rect 162766 7982 162818 8034
rect 162818 7982 162820 8034
rect 162764 7980 162820 7982
rect 163548 11116 163604 11172
rect 163772 11004 163828 11060
rect 163996 10780 164052 10836
rect 164444 10834 164500 10836
rect 164444 10782 164446 10834
rect 164446 10782 164498 10834
rect 164498 10782 164500 10834
rect 164444 10780 164500 10782
rect 168028 14364 168084 14420
rect 173436 45498 173492 45500
rect 173436 45446 173438 45498
rect 173438 45446 173490 45498
rect 173490 45446 173492 45498
rect 173436 45444 173492 45446
rect 173540 45498 173596 45500
rect 173540 45446 173542 45498
rect 173542 45446 173594 45498
rect 173594 45446 173596 45498
rect 173540 45444 173596 45446
rect 173644 45498 173700 45500
rect 173644 45446 173646 45498
rect 173646 45446 173698 45498
rect 173698 45446 173700 45498
rect 173644 45444 173700 45446
rect 173436 43930 173492 43932
rect 173436 43878 173438 43930
rect 173438 43878 173490 43930
rect 173490 43878 173492 43930
rect 173436 43876 173492 43878
rect 173540 43930 173596 43932
rect 173540 43878 173542 43930
rect 173542 43878 173594 43930
rect 173594 43878 173596 43930
rect 173540 43876 173596 43878
rect 173644 43930 173700 43932
rect 173644 43878 173646 43930
rect 173646 43878 173698 43930
rect 173698 43878 173700 43930
rect 173644 43876 173700 43878
rect 173068 43708 173124 43764
rect 173436 42362 173492 42364
rect 173436 42310 173438 42362
rect 173438 42310 173490 42362
rect 173490 42310 173492 42362
rect 173436 42308 173492 42310
rect 173540 42362 173596 42364
rect 173540 42310 173542 42362
rect 173542 42310 173594 42362
rect 173594 42310 173596 42362
rect 173540 42308 173596 42310
rect 173644 42362 173700 42364
rect 173644 42310 173646 42362
rect 173646 42310 173698 42362
rect 173698 42310 173700 42362
rect 173644 42308 173700 42310
rect 173436 40794 173492 40796
rect 173436 40742 173438 40794
rect 173438 40742 173490 40794
rect 173490 40742 173492 40794
rect 173436 40740 173492 40742
rect 173540 40794 173596 40796
rect 173540 40742 173542 40794
rect 173542 40742 173594 40794
rect 173594 40742 173596 40794
rect 173540 40740 173596 40742
rect 173644 40794 173700 40796
rect 173644 40742 173646 40794
rect 173646 40742 173698 40794
rect 173698 40742 173700 40794
rect 173644 40740 173700 40742
rect 173436 39226 173492 39228
rect 173436 39174 173438 39226
rect 173438 39174 173490 39226
rect 173490 39174 173492 39226
rect 173436 39172 173492 39174
rect 173540 39226 173596 39228
rect 173540 39174 173542 39226
rect 173542 39174 173594 39226
rect 173594 39174 173596 39226
rect 173540 39172 173596 39174
rect 173644 39226 173700 39228
rect 173644 39174 173646 39226
rect 173646 39174 173698 39226
rect 173698 39174 173700 39226
rect 173644 39172 173700 39174
rect 173436 37658 173492 37660
rect 173436 37606 173438 37658
rect 173438 37606 173490 37658
rect 173490 37606 173492 37658
rect 173436 37604 173492 37606
rect 173540 37658 173596 37660
rect 173540 37606 173542 37658
rect 173542 37606 173594 37658
rect 173594 37606 173596 37658
rect 173540 37604 173596 37606
rect 173644 37658 173700 37660
rect 173644 37606 173646 37658
rect 173646 37606 173698 37658
rect 173698 37606 173700 37658
rect 173644 37604 173700 37606
rect 173436 36090 173492 36092
rect 173436 36038 173438 36090
rect 173438 36038 173490 36090
rect 173490 36038 173492 36090
rect 173436 36036 173492 36038
rect 173540 36090 173596 36092
rect 173540 36038 173542 36090
rect 173542 36038 173594 36090
rect 173594 36038 173596 36090
rect 173540 36036 173596 36038
rect 173644 36090 173700 36092
rect 173644 36038 173646 36090
rect 173646 36038 173698 36090
rect 173698 36038 173700 36090
rect 173644 36036 173700 36038
rect 173436 34522 173492 34524
rect 173436 34470 173438 34522
rect 173438 34470 173490 34522
rect 173490 34470 173492 34522
rect 173436 34468 173492 34470
rect 173540 34522 173596 34524
rect 173540 34470 173542 34522
rect 173542 34470 173594 34522
rect 173594 34470 173596 34522
rect 173540 34468 173596 34470
rect 173644 34522 173700 34524
rect 173644 34470 173646 34522
rect 173646 34470 173698 34522
rect 173698 34470 173700 34522
rect 173644 34468 173700 34470
rect 173436 32954 173492 32956
rect 173436 32902 173438 32954
rect 173438 32902 173490 32954
rect 173490 32902 173492 32954
rect 173436 32900 173492 32902
rect 173540 32954 173596 32956
rect 173540 32902 173542 32954
rect 173542 32902 173594 32954
rect 173594 32902 173596 32954
rect 173540 32900 173596 32902
rect 173644 32954 173700 32956
rect 173644 32902 173646 32954
rect 173646 32902 173698 32954
rect 173698 32902 173700 32954
rect 173644 32900 173700 32902
rect 173436 31386 173492 31388
rect 173436 31334 173438 31386
rect 173438 31334 173490 31386
rect 173490 31334 173492 31386
rect 173436 31332 173492 31334
rect 173540 31386 173596 31388
rect 173540 31334 173542 31386
rect 173542 31334 173594 31386
rect 173594 31334 173596 31386
rect 173540 31332 173596 31334
rect 173644 31386 173700 31388
rect 173644 31334 173646 31386
rect 173646 31334 173698 31386
rect 173698 31334 173700 31386
rect 173644 31332 173700 31334
rect 173436 29818 173492 29820
rect 173436 29766 173438 29818
rect 173438 29766 173490 29818
rect 173490 29766 173492 29818
rect 173436 29764 173492 29766
rect 173540 29818 173596 29820
rect 173540 29766 173542 29818
rect 173542 29766 173594 29818
rect 173594 29766 173596 29818
rect 173540 29764 173596 29766
rect 173644 29818 173700 29820
rect 173644 29766 173646 29818
rect 173646 29766 173698 29818
rect 173698 29766 173700 29818
rect 173644 29764 173700 29766
rect 173436 28250 173492 28252
rect 173436 28198 173438 28250
rect 173438 28198 173490 28250
rect 173490 28198 173492 28250
rect 173436 28196 173492 28198
rect 173540 28250 173596 28252
rect 173540 28198 173542 28250
rect 173542 28198 173594 28250
rect 173594 28198 173596 28250
rect 173540 28196 173596 28198
rect 173644 28250 173700 28252
rect 173644 28198 173646 28250
rect 173646 28198 173698 28250
rect 173698 28198 173700 28250
rect 173644 28196 173700 28198
rect 173436 26682 173492 26684
rect 173436 26630 173438 26682
rect 173438 26630 173490 26682
rect 173490 26630 173492 26682
rect 173436 26628 173492 26630
rect 173540 26682 173596 26684
rect 173540 26630 173542 26682
rect 173542 26630 173594 26682
rect 173594 26630 173596 26682
rect 173540 26628 173596 26630
rect 173644 26682 173700 26684
rect 173644 26630 173646 26682
rect 173646 26630 173698 26682
rect 173698 26630 173700 26682
rect 173644 26628 173700 26630
rect 173436 25114 173492 25116
rect 173436 25062 173438 25114
rect 173438 25062 173490 25114
rect 173490 25062 173492 25114
rect 173436 25060 173492 25062
rect 173540 25114 173596 25116
rect 173540 25062 173542 25114
rect 173542 25062 173594 25114
rect 173594 25062 173596 25114
rect 173540 25060 173596 25062
rect 173644 25114 173700 25116
rect 173644 25062 173646 25114
rect 173646 25062 173698 25114
rect 173698 25062 173700 25114
rect 173644 25060 173700 25062
rect 173436 23546 173492 23548
rect 173436 23494 173438 23546
rect 173438 23494 173490 23546
rect 173490 23494 173492 23546
rect 173436 23492 173492 23494
rect 173540 23546 173596 23548
rect 173540 23494 173542 23546
rect 173542 23494 173594 23546
rect 173594 23494 173596 23546
rect 173540 23492 173596 23494
rect 173644 23546 173700 23548
rect 173644 23494 173646 23546
rect 173646 23494 173698 23546
rect 173698 23494 173700 23546
rect 173644 23492 173700 23494
rect 173436 21978 173492 21980
rect 173436 21926 173438 21978
rect 173438 21926 173490 21978
rect 173490 21926 173492 21978
rect 173436 21924 173492 21926
rect 173540 21978 173596 21980
rect 173540 21926 173542 21978
rect 173542 21926 173594 21978
rect 173594 21926 173596 21978
rect 173540 21924 173596 21926
rect 173644 21978 173700 21980
rect 173644 21926 173646 21978
rect 173646 21926 173698 21978
rect 173698 21926 173700 21978
rect 173644 21924 173700 21926
rect 173436 20410 173492 20412
rect 173436 20358 173438 20410
rect 173438 20358 173490 20410
rect 173490 20358 173492 20410
rect 173436 20356 173492 20358
rect 173540 20410 173596 20412
rect 173540 20358 173542 20410
rect 173542 20358 173594 20410
rect 173594 20358 173596 20410
rect 173540 20356 173596 20358
rect 173644 20410 173700 20412
rect 173644 20358 173646 20410
rect 173646 20358 173698 20410
rect 173698 20358 173700 20410
rect 173644 20356 173700 20358
rect 173436 18842 173492 18844
rect 173436 18790 173438 18842
rect 173438 18790 173490 18842
rect 173490 18790 173492 18842
rect 173436 18788 173492 18790
rect 173540 18842 173596 18844
rect 173540 18790 173542 18842
rect 173542 18790 173594 18842
rect 173594 18790 173596 18842
rect 173540 18788 173596 18790
rect 173644 18842 173700 18844
rect 173644 18790 173646 18842
rect 173646 18790 173698 18842
rect 173698 18790 173700 18842
rect 173644 18788 173700 18790
rect 173436 17274 173492 17276
rect 173436 17222 173438 17274
rect 173438 17222 173490 17274
rect 173490 17222 173492 17274
rect 173436 17220 173492 17222
rect 173540 17274 173596 17276
rect 173540 17222 173542 17274
rect 173542 17222 173594 17274
rect 173594 17222 173596 17274
rect 173540 17220 173596 17222
rect 173644 17274 173700 17276
rect 173644 17222 173646 17274
rect 173646 17222 173698 17274
rect 173698 17222 173700 17274
rect 173644 17220 173700 17222
rect 173436 15706 173492 15708
rect 173436 15654 173438 15706
rect 173438 15654 173490 15706
rect 173490 15654 173492 15706
rect 173436 15652 173492 15654
rect 173540 15706 173596 15708
rect 173540 15654 173542 15706
rect 173542 15654 173594 15706
rect 173594 15654 173596 15706
rect 173540 15652 173596 15654
rect 173644 15706 173700 15708
rect 173644 15654 173646 15706
rect 173646 15654 173698 15706
rect 173698 15654 173700 15706
rect 173644 15652 173700 15654
rect 169260 14140 169316 14196
rect 173436 14138 173492 14140
rect 173436 14086 173438 14138
rect 173438 14086 173490 14138
rect 173490 14086 173492 14138
rect 173436 14084 173492 14086
rect 173540 14138 173596 14140
rect 173540 14086 173542 14138
rect 173542 14086 173594 14138
rect 173594 14086 173596 14138
rect 173540 14084 173596 14086
rect 173644 14138 173700 14140
rect 173644 14086 173646 14138
rect 173646 14086 173698 14138
rect 173698 14086 173700 14138
rect 173644 14084 173700 14086
rect 173436 12570 173492 12572
rect 173436 12518 173438 12570
rect 173438 12518 173490 12570
rect 173490 12518 173492 12570
rect 173436 12516 173492 12518
rect 173540 12570 173596 12572
rect 173540 12518 173542 12570
rect 173542 12518 173594 12570
rect 173594 12518 173596 12570
rect 173540 12516 173596 12518
rect 173644 12570 173700 12572
rect 173644 12518 173646 12570
rect 173646 12518 173698 12570
rect 173698 12518 173700 12570
rect 173644 12516 173700 12518
rect 180684 14364 180740 14420
rect 182252 45500 182308 45556
rect 176876 12012 176932 12068
rect 168028 11676 168084 11732
rect 173436 11002 173492 11004
rect 173436 10950 173438 11002
rect 173438 10950 173490 11002
rect 173490 10950 173492 11002
rect 173436 10948 173492 10950
rect 173540 11002 173596 11004
rect 173540 10950 173542 11002
rect 173542 10950 173594 11002
rect 173594 10950 173596 11002
rect 173540 10948 173596 10950
rect 173644 11002 173700 11004
rect 173644 10950 173646 11002
rect 173646 10950 173698 11002
rect 173698 10950 173700 11002
rect 173644 10948 173700 10950
rect 167132 10780 167188 10836
rect 163324 10610 163380 10612
rect 163324 10558 163326 10610
rect 163326 10558 163378 10610
rect 163378 10558 163380 10610
rect 163324 10556 163380 10558
rect 173436 9434 173492 9436
rect 173436 9382 173438 9434
rect 173438 9382 173490 9434
rect 173490 9382 173492 9434
rect 173436 9380 173492 9382
rect 173540 9434 173596 9436
rect 173540 9382 173542 9434
rect 173542 9382 173594 9434
rect 173594 9382 173596 9434
rect 173540 9380 173596 9382
rect 173644 9434 173700 9436
rect 173644 9382 173646 9434
rect 173646 9382 173698 9434
rect 173698 9382 173700 9434
rect 173644 9380 173700 9382
rect 163436 8428 163492 8484
rect 163996 8540 164052 8596
rect 162652 7084 162708 7140
rect 162428 6972 162484 7028
rect 162988 7532 163044 7588
rect 162764 6972 162820 7028
rect 162652 6690 162708 6692
rect 162652 6638 162654 6690
rect 162654 6638 162706 6690
rect 162706 6638 162708 6690
rect 162652 6636 162708 6638
rect 162876 6578 162932 6580
rect 162876 6526 162878 6578
rect 162878 6526 162930 6578
rect 162930 6526 162932 6578
rect 162876 6524 162932 6526
rect 162764 6076 162820 6132
rect 162316 5404 162372 5460
rect 163100 6524 163156 6580
rect 162876 5292 162932 5348
rect 163324 6748 163380 6804
rect 163324 6188 163380 6244
rect 163100 5292 163156 5348
rect 162988 5010 163044 5012
rect 162988 4958 162990 5010
rect 162990 4958 163042 5010
rect 163042 4958 163044 5010
rect 162988 4956 163044 4958
rect 163324 5180 163380 5236
rect 161980 4620 162036 4676
rect 162204 4396 162260 4452
rect 162764 4450 162820 4452
rect 162764 4398 162766 4450
rect 162766 4398 162818 4450
rect 162818 4398 162820 4450
rect 162764 4396 162820 4398
rect 163548 6076 163604 6132
rect 163548 5404 163604 5460
rect 163884 6524 163940 6580
rect 163772 6466 163828 6468
rect 163772 6414 163774 6466
rect 163774 6414 163826 6466
rect 163826 6414 163828 6466
rect 163772 6412 163828 6414
rect 164332 7980 164388 8036
rect 163996 6412 164052 6468
rect 164220 6636 164276 6692
rect 173436 7866 173492 7868
rect 173436 7814 173438 7866
rect 173438 7814 173490 7866
rect 173490 7814 173492 7866
rect 173436 7812 173492 7814
rect 173540 7866 173596 7868
rect 173540 7814 173542 7866
rect 173542 7814 173594 7866
rect 173594 7814 173596 7866
rect 173540 7812 173596 7814
rect 173644 7866 173700 7868
rect 173644 7814 173646 7866
rect 173646 7814 173698 7866
rect 173698 7814 173700 7866
rect 173644 7812 173700 7814
rect 170492 7308 170548 7364
rect 167804 6748 167860 6804
rect 164556 6466 164612 6468
rect 164556 6414 164558 6466
rect 164558 6414 164610 6466
rect 164610 6414 164612 6466
rect 164556 6412 164612 6414
rect 164220 6076 164276 6132
rect 163996 6018 164052 6020
rect 163996 5966 163998 6018
rect 163998 5966 164050 6018
rect 164050 5966 164052 6018
rect 163996 5964 164052 5966
rect 164108 5906 164164 5908
rect 164108 5854 164110 5906
rect 164110 5854 164162 5906
rect 164162 5854 164164 5906
rect 164108 5852 164164 5854
rect 163772 5740 163828 5796
rect 163772 5516 163828 5572
rect 163996 5180 164052 5236
rect 163772 4844 163828 4900
rect 163660 4562 163716 4564
rect 163660 4510 163662 4562
rect 163662 4510 163714 4562
rect 163714 4510 163716 4562
rect 163660 4508 163716 4510
rect 164220 4620 164276 4676
rect 163996 4338 164052 4340
rect 163996 4286 163998 4338
rect 163998 4286 164050 4338
rect 164050 4286 164052 4338
rect 163996 4284 164052 4286
rect 161644 3836 161700 3892
rect 161980 3442 162036 3444
rect 161980 3390 161982 3442
rect 161982 3390 162034 3442
rect 162034 3390 162036 3442
rect 161980 3388 162036 3390
rect 160748 2716 160804 2772
rect 163324 3836 163380 3892
rect 164556 5516 164612 5572
rect 165116 6466 165172 6468
rect 165116 6414 165118 6466
rect 165118 6414 165170 6466
rect 165170 6414 165172 6466
rect 165116 6412 165172 6414
rect 164444 5404 164500 5460
rect 164780 5292 164836 5348
rect 165116 5906 165172 5908
rect 165116 5854 165118 5906
rect 165118 5854 165170 5906
rect 165170 5854 165172 5906
rect 165116 5852 165172 5854
rect 165564 5906 165620 5908
rect 165564 5854 165566 5906
rect 165566 5854 165618 5906
rect 165618 5854 165620 5906
rect 165564 5852 165620 5854
rect 165004 5628 165060 5684
rect 165676 5292 165732 5348
rect 165228 5180 165284 5236
rect 166124 5180 166180 5236
rect 166236 5122 166292 5124
rect 166236 5070 166238 5122
rect 166238 5070 166290 5122
rect 166290 5070 166292 5122
rect 166236 5068 166292 5070
rect 164332 3836 164388 3892
rect 163660 3442 163716 3444
rect 163660 3390 163662 3442
rect 163662 3390 163714 3442
rect 163714 3390 163716 3442
rect 163660 3388 163716 3390
rect 163212 2940 163268 2996
rect 165340 4396 165396 4452
rect 165452 4284 165508 4340
rect 165676 4226 165732 4228
rect 165676 4174 165678 4226
rect 165678 4174 165730 4226
rect 165730 4174 165732 4226
rect 165676 4172 165732 4174
rect 166908 3612 166964 3668
rect 164444 2828 164500 2884
rect 167580 3442 167636 3444
rect 167580 3390 167582 3442
rect 167582 3390 167634 3442
rect 167634 3390 167636 3442
rect 167580 3388 167636 3390
rect 168140 3442 168196 3444
rect 168140 3390 168142 3442
rect 168142 3390 168194 3442
rect 168194 3390 168196 3442
rect 168140 3388 168196 3390
rect 173436 6298 173492 6300
rect 173436 6246 173438 6298
rect 173438 6246 173490 6298
rect 173490 6246 173492 6298
rect 173436 6244 173492 6246
rect 173540 6298 173596 6300
rect 173540 6246 173542 6298
rect 173542 6246 173594 6298
rect 173594 6246 173596 6298
rect 173540 6244 173596 6246
rect 173644 6298 173700 6300
rect 173644 6246 173646 6298
rect 173646 6246 173698 6298
rect 173698 6246 173700 6298
rect 173644 6244 173700 6246
rect 181244 5852 181300 5908
rect 178556 4956 178612 5012
rect 173436 4730 173492 4732
rect 173436 4678 173438 4730
rect 173438 4678 173490 4730
rect 173490 4678 173492 4730
rect 173436 4676 173492 4678
rect 173540 4730 173596 4732
rect 173540 4678 173542 4730
rect 173542 4678 173594 4730
rect 173594 4678 173596 4730
rect 173540 4676 173596 4678
rect 173644 4730 173700 4732
rect 173644 4678 173646 4730
rect 173646 4678 173698 4730
rect 173698 4678 173700 4730
rect 173644 4676 173700 4678
rect 175868 3836 175924 3892
rect 173180 3724 173236 3780
rect 172956 3388 173012 3444
rect 173516 3442 173572 3444
rect 173516 3390 173518 3442
rect 173518 3390 173570 3442
rect 173570 3390 173572 3442
rect 173516 3388 173572 3390
rect 173436 3162 173492 3164
rect 173436 3110 173438 3162
rect 173438 3110 173490 3162
rect 173490 3110 173492 3162
rect 173436 3108 173492 3110
rect 173540 3162 173596 3164
rect 173540 3110 173542 3162
rect 173542 3110 173594 3162
rect 173594 3110 173596 3162
rect 173540 3108 173596 3110
rect 173644 3162 173700 3164
rect 173644 3110 173646 3162
rect 173646 3110 173698 3162
rect 173698 3110 173700 3162
rect 173644 3108 173700 3110
rect 181020 3442 181076 3444
rect 181020 3390 181022 3442
rect 181022 3390 181074 3442
rect 181074 3390 181076 3442
rect 181020 3388 181076 3390
rect 181580 3442 181636 3444
rect 181580 3390 181582 3442
rect 181582 3390 181634 3442
rect 181634 3390 181636 3442
rect 181580 3388 181636 3390
rect 184604 15932 184660 15988
rect 189196 45778 189252 45780
rect 189196 45726 189198 45778
rect 189198 45726 189250 45778
rect 189250 45726 189252 45778
rect 189196 45724 189252 45726
rect 188796 44714 188852 44716
rect 188796 44662 188798 44714
rect 188798 44662 188850 44714
rect 188850 44662 188852 44714
rect 188796 44660 188852 44662
rect 188900 44714 188956 44716
rect 188900 44662 188902 44714
rect 188902 44662 188954 44714
rect 188954 44662 188956 44714
rect 188900 44660 188956 44662
rect 189004 44714 189060 44716
rect 189004 44662 189006 44714
rect 189006 44662 189058 44714
rect 189058 44662 189060 44714
rect 189004 44660 189060 44662
rect 188796 43146 188852 43148
rect 188796 43094 188798 43146
rect 188798 43094 188850 43146
rect 188850 43094 188852 43146
rect 188796 43092 188852 43094
rect 188900 43146 188956 43148
rect 188900 43094 188902 43146
rect 188902 43094 188954 43146
rect 188954 43094 188956 43146
rect 188900 43092 188956 43094
rect 189004 43146 189060 43148
rect 189004 43094 189006 43146
rect 189006 43094 189058 43146
rect 189058 43094 189060 43146
rect 189004 43092 189060 43094
rect 188796 41578 188852 41580
rect 188796 41526 188798 41578
rect 188798 41526 188850 41578
rect 188850 41526 188852 41578
rect 188796 41524 188852 41526
rect 188900 41578 188956 41580
rect 188900 41526 188902 41578
rect 188902 41526 188954 41578
rect 188954 41526 188956 41578
rect 188900 41524 188956 41526
rect 189004 41578 189060 41580
rect 189004 41526 189006 41578
rect 189006 41526 189058 41578
rect 189058 41526 189060 41578
rect 189004 41524 189060 41526
rect 188796 40010 188852 40012
rect 188796 39958 188798 40010
rect 188798 39958 188850 40010
rect 188850 39958 188852 40010
rect 188796 39956 188852 39958
rect 188900 40010 188956 40012
rect 188900 39958 188902 40010
rect 188902 39958 188954 40010
rect 188954 39958 188956 40010
rect 188900 39956 188956 39958
rect 189004 40010 189060 40012
rect 189004 39958 189006 40010
rect 189006 39958 189058 40010
rect 189058 39958 189060 40010
rect 189004 39956 189060 39958
rect 188796 38442 188852 38444
rect 188796 38390 188798 38442
rect 188798 38390 188850 38442
rect 188850 38390 188852 38442
rect 188796 38388 188852 38390
rect 188900 38442 188956 38444
rect 188900 38390 188902 38442
rect 188902 38390 188954 38442
rect 188954 38390 188956 38442
rect 188900 38388 188956 38390
rect 189004 38442 189060 38444
rect 189004 38390 189006 38442
rect 189006 38390 189058 38442
rect 189058 38390 189060 38442
rect 189004 38388 189060 38390
rect 188796 36874 188852 36876
rect 188796 36822 188798 36874
rect 188798 36822 188850 36874
rect 188850 36822 188852 36874
rect 188796 36820 188852 36822
rect 188900 36874 188956 36876
rect 188900 36822 188902 36874
rect 188902 36822 188954 36874
rect 188954 36822 188956 36874
rect 188900 36820 188956 36822
rect 189004 36874 189060 36876
rect 189004 36822 189006 36874
rect 189006 36822 189058 36874
rect 189058 36822 189060 36874
rect 189004 36820 189060 36822
rect 188796 35306 188852 35308
rect 188796 35254 188798 35306
rect 188798 35254 188850 35306
rect 188850 35254 188852 35306
rect 188796 35252 188852 35254
rect 188900 35306 188956 35308
rect 188900 35254 188902 35306
rect 188902 35254 188954 35306
rect 188954 35254 188956 35306
rect 188900 35252 188956 35254
rect 189004 35306 189060 35308
rect 189004 35254 189006 35306
rect 189006 35254 189058 35306
rect 189058 35254 189060 35306
rect 189004 35252 189060 35254
rect 188796 33738 188852 33740
rect 188796 33686 188798 33738
rect 188798 33686 188850 33738
rect 188850 33686 188852 33738
rect 188796 33684 188852 33686
rect 188900 33738 188956 33740
rect 188900 33686 188902 33738
rect 188902 33686 188954 33738
rect 188954 33686 188956 33738
rect 188900 33684 188956 33686
rect 189004 33738 189060 33740
rect 189004 33686 189006 33738
rect 189006 33686 189058 33738
rect 189058 33686 189060 33738
rect 189004 33684 189060 33686
rect 188796 32170 188852 32172
rect 188796 32118 188798 32170
rect 188798 32118 188850 32170
rect 188850 32118 188852 32170
rect 188796 32116 188852 32118
rect 188900 32170 188956 32172
rect 188900 32118 188902 32170
rect 188902 32118 188954 32170
rect 188954 32118 188956 32170
rect 188900 32116 188956 32118
rect 189004 32170 189060 32172
rect 189004 32118 189006 32170
rect 189006 32118 189058 32170
rect 189058 32118 189060 32170
rect 189004 32116 189060 32118
rect 188796 30602 188852 30604
rect 188796 30550 188798 30602
rect 188798 30550 188850 30602
rect 188850 30550 188852 30602
rect 188796 30548 188852 30550
rect 188900 30602 188956 30604
rect 188900 30550 188902 30602
rect 188902 30550 188954 30602
rect 188954 30550 188956 30602
rect 188900 30548 188956 30550
rect 189004 30602 189060 30604
rect 189004 30550 189006 30602
rect 189006 30550 189058 30602
rect 189058 30550 189060 30602
rect 189004 30548 189060 30550
rect 188796 29034 188852 29036
rect 188796 28982 188798 29034
rect 188798 28982 188850 29034
rect 188850 28982 188852 29034
rect 188796 28980 188852 28982
rect 188900 29034 188956 29036
rect 188900 28982 188902 29034
rect 188902 28982 188954 29034
rect 188954 28982 188956 29034
rect 188900 28980 188956 28982
rect 189004 29034 189060 29036
rect 189004 28982 189006 29034
rect 189006 28982 189058 29034
rect 189058 28982 189060 29034
rect 189004 28980 189060 28982
rect 188796 27466 188852 27468
rect 188796 27414 188798 27466
rect 188798 27414 188850 27466
rect 188850 27414 188852 27466
rect 188796 27412 188852 27414
rect 188900 27466 188956 27468
rect 188900 27414 188902 27466
rect 188902 27414 188954 27466
rect 188954 27414 188956 27466
rect 188900 27412 188956 27414
rect 189004 27466 189060 27468
rect 189004 27414 189006 27466
rect 189006 27414 189058 27466
rect 189058 27414 189060 27466
rect 189004 27412 189060 27414
rect 188796 25898 188852 25900
rect 188796 25846 188798 25898
rect 188798 25846 188850 25898
rect 188850 25846 188852 25898
rect 188796 25844 188852 25846
rect 188900 25898 188956 25900
rect 188900 25846 188902 25898
rect 188902 25846 188954 25898
rect 188954 25846 188956 25898
rect 188900 25844 188956 25846
rect 189004 25898 189060 25900
rect 189004 25846 189006 25898
rect 189006 25846 189058 25898
rect 189058 25846 189060 25898
rect 189004 25844 189060 25846
rect 188796 24330 188852 24332
rect 188796 24278 188798 24330
rect 188798 24278 188850 24330
rect 188850 24278 188852 24330
rect 188796 24276 188852 24278
rect 188900 24330 188956 24332
rect 188900 24278 188902 24330
rect 188902 24278 188954 24330
rect 188954 24278 188956 24330
rect 188900 24276 188956 24278
rect 189004 24330 189060 24332
rect 189004 24278 189006 24330
rect 189006 24278 189058 24330
rect 189058 24278 189060 24330
rect 189004 24276 189060 24278
rect 188796 22762 188852 22764
rect 188796 22710 188798 22762
rect 188798 22710 188850 22762
rect 188850 22710 188852 22762
rect 188796 22708 188852 22710
rect 188900 22762 188956 22764
rect 188900 22710 188902 22762
rect 188902 22710 188954 22762
rect 188954 22710 188956 22762
rect 188900 22708 188956 22710
rect 189004 22762 189060 22764
rect 189004 22710 189006 22762
rect 189006 22710 189058 22762
rect 189058 22710 189060 22762
rect 189004 22708 189060 22710
rect 188796 21194 188852 21196
rect 188796 21142 188798 21194
rect 188798 21142 188850 21194
rect 188850 21142 188852 21194
rect 188796 21140 188852 21142
rect 188900 21194 188956 21196
rect 188900 21142 188902 21194
rect 188902 21142 188954 21194
rect 188954 21142 188956 21194
rect 188900 21140 188956 21142
rect 189004 21194 189060 21196
rect 189004 21142 189006 21194
rect 189006 21142 189058 21194
rect 189058 21142 189060 21194
rect 189004 21140 189060 21142
rect 188796 19626 188852 19628
rect 188796 19574 188798 19626
rect 188798 19574 188850 19626
rect 188850 19574 188852 19626
rect 188796 19572 188852 19574
rect 188900 19626 188956 19628
rect 188900 19574 188902 19626
rect 188902 19574 188954 19626
rect 188954 19574 188956 19626
rect 188900 19572 188956 19574
rect 189004 19626 189060 19628
rect 189004 19574 189006 19626
rect 189006 19574 189058 19626
rect 189058 19574 189060 19626
rect 189004 19572 189060 19574
rect 188796 18058 188852 18060
rect 188796 18006 188798 18058
rect 188798 18006 188850 18058
rect 188850 18006 188852 18058
rect 188796 18004 188852 18006
rect 188900 18058 188956 18060
rect 188900 18006 188902 18058
rect 188902 18006 188954 18058
rect 188954 18006 188956 18058
rect 188900 18004 188956 18006
rect 189004 18058 189060 18060
rect 189004 18006 189006 18058
rect 189006 18006 189058 18058
rect 189058 18006 189060 18058
rect 189004 18004 189060 18006
rect 188796 16490 188852 16492
rect 188796 16438 188798 16490
rect 188798 16438 188850 16490
rect 188850 16438 188852 16490
rect 188796 16436 188852 16438
rect 188900 16490 188956 16492
rect 188900 16438 188902 16490
rect 188902 16438 188954 16490
rect 188954 16438 188956 16490
rect 188900 16436 188956 16438
rect 189004 16490 189060 16492
rect 189004 16438 189006 16490
rect 189006 16438 189058 16490
rect 189058 16438 189060 16490
rect 189004 16436 189060 16438
rect 188796 14922 188852 14924
rect 188796 14870 188798 14922
rect 188798 14870 188850 14922
rect 188850 14870 188852 14922
rect 188796 14868 188852 14870
rect 188900 14922 188956 14924
rect 188900 14870 188902 14922
rect 188902 14870 188954 14922
rect 188954 14870 188956 14922
rect 188900 14868 188956 14870
rect 189004 14922 189060 14924
rect 189004 14870 189006 14922
rect 189006 14870 189058 14922
rect 189058 14870 189060 14922
rect 189004 14868 189060 14870
rect 188796 13354 188852 13356
rect 188796 13302 188798 13354
rect 188798 13302 188850 13354
rect 188850 13302 188852 13354
rect 188796 13300 188852 13302
rect 188900 13354 188956 13356
rect 188900 13302 188902 13354
rect 188902 13302 188954 13354
rect 188954 13302 188956 13354
rect 188900 13300 188956 13302
rect 189004 13354 189060 13356
rect 189004 13302 189006 13354
rect 189006 13302 189058 13354
rect 189058 13302 189060 13354
rect 189004 13300 189060 13302
rect 187292 12908 187348 12964
rect 205212 46002 205268 46004
rect 205212 45950 205214 46002
rect 205214 45950 205266 46002
rect 205266 45950 205268 46002
rect 205212 45948 205268 45950
rect 205772 45948 205828 46004
rect 201292 45778 201348 45780
rect 201292 45726 201294 45778
rect 201294 45726 201346 45778
rect 201346 45726 201348 45778
rect 201292 45724 201348 45726
rect 204156 45498 204212 45500
rect 204156 45446 204158 45498
rect 204158 45446 204210 45498
rect 204210 45446 204212 45498
rect 204156 45444 204212 45446
rect 204260 45498 204316 45500
rect 204260 45446 204262 45498
rect 204262 45446 204314 45498
rect 204314 45446 204316 45498
rect 204260 45444 204316 45446
rect 204364 45498 204420 45500
rect 204364 45446 204366 45498
rect 204366 45446 204418 45498
rect 204418 45446 204420 45498
rect 204364 45444 204420 45446
rect 204156 43930 204212 43932
rect 204156 43878 204158 43930
rect 204158 43878 204210 43930
rect 204210 43878 204212 43930
rect 204156 43876 204212 43878
rect 204260 43930 204316 43932
rect 204260 43878 204262 43930
rect 204262 43878 204314 43930
rect 204314 43878 204316 43930
rect 204260 43876 204316 43878
rect 204364 43930 204420 43932
rect 204364 43878 204366 43930
rect 204366 43878 204418 43930
rect 204418 43878 204420 43930
rect 204364 43876 204420 43878
rect 204156 42362 204212 42364
rect 204156 42310 204158 42362
rect 204158 42310 204210 42362
rect 204210 42310 204212 42362
rect 204156 42308 204212 42310
rect 204260 42362 204316 42364
rect 204260 42310 204262 42362
rect 204262 42310 204314 42362
rect 204314 42310 204316 42362
rect 204260 42308 204316 42310
rect 204364 42362 204420 42364
rect 204364 42310 204366 42362
rect 204366 42310 204418 42362
rect 204418 42310 204420 42362
rect 204364 42308 204420 42310
rect 204156 40794 204212 40796
rect 204156 40742 204158 40794
rect 204158 40742 204210 40794
rect 204210 40742 204212 40794
rect 204156 40740 204212 40742
rect 204260 40794 204316 40796
rect 204260 40742 204262 40794
rect 204262 40742 204314 40794
rect 204314 40742 204316 40794
rect 204260 40740 204316 40742
rect 204364 40794 204420 40796
rect 204364 40742 204366 40794
rect 204366 40742 204418 40794
rect 204418 40742 204420 40794
rect 204364 40740 204420 40742
rect 204156 39226 204212 39228
rect 204156 39174 204158 39226
rect 204158 39174 204210 39226
rect 204210 39174 204212 39226
rect 204156 39172 204212 39174
rect 204260 39226 204316 39228
rect 204260 39174 204262 39226
rect 204262 39174 204314 39226
rect 204314 39174 204316 39226
rect 204260 39172 204316 39174
rect 204364 39226 204420 39228
rect 204364 39174 204366 39226
rect 204366 39174 204418 39226
rect 204418 39174 204420 39226
rect 204364 39172 204420 39174
rect 204156 37658 204212 37660
rect 204156 37606 204158 37658
rect 204158 37606 204210 37658
rect 204210 37606 204212 37658
rect 204156 37604 204212 37606
rect 204260 37658 204316 37660
rect 204260 37606 204262 37658
rect 204262 37606 204314 37658
rect 204314 37606 204316 37658
rect 204260 37604 204316 37606
rect 204364 37658 204420 37660
rect 204364 37606 204366 37658
rect 204366 37606 204418 37658
rect 204418 37606 204420 37658
rect 204364 37604 204420 37606
rect 204156 36090 204212 36092
rect 204156 36038 204158 36090
rect 204158 36038 204210 36090
rect 204210 36038 204212 36090
rect 204156 36036 204212 36038
rect 204260 36090 204316 36092
rect 204260 36038 204262 36090
rect 204262 36038 204314 36090
rect 204314 36038 204316 36090
rect 204260 36036 204316 36038
rect 204364 36090 204420 36092
rect 204364 36038 204366 36090
rect 204366 36038 204418 36090
rect 204418 36038 204420 36090
rect 204364 36036 204420 36038
rect 204156 34522 204212 34524
rect 204156 34470 204158 34522
rect 204158 34470 204210 34522
rect 204210 34470 204212 34522
rect 204156 34468 204212 34470
rect 204260 34522 204316 34524
rect 204260 34470 204262 34522
rect 204262 34470 204314 34522
rect 204314 34470 204316 34522
rect 204260 34468 204316 34470
rect 204364 34522 204420 34524
rect 204364 34470 204366 34522
rect 204366 34470 204418 34522
rect 204418 34470 204420 34522
rect 204364 34468 204420 34470
rect 204156 32954 204212 32956
rect 204156 32902 204158 32954
rect 204158 32902 204210 32954
rect 204210 32902 204212 32954
rect 204156 32900 204212 32902
rect 204260 32954 204316 32956
rect 204260 32902 204262 32954
rect 204262 32902 204314 32954
rect 204314 32902 204316 32954
rect 204260 32900 204316 32902
rect 204364 32954 204420 32956
rect 204364 32902 204366 32954
rect 204366 32902 204418 32954
rect 204418 32902 204420 32954
rect 204364 32900 204420 32902
rect 204156 31386 204212 31388
rect 204156 31334 204158 31386
rect 204158 31334 204210 31386
rect 204210 31334 204212 31386
rect 204156 31332 204212 31334
rect 204260 31386 204316 31388
rect 204260 31334 204262 31386
rect 204262 31334 204314 31386
rect 204314 31334 204316 31386
rect 204260 31332 204316 31334
rect 204364 31386 204420 31388
rect 204364 31334 204366 31386
rect 204366 31334 204418 31386
rect 204418 31334 204420 31386
rect 204364 31332 204420 31334
rect 204156 29818 204212 29820
rect 204156 29766 204158 29818
rect 204158 29766 204210 29818
rect 204210 29766 204212 29818
rect 204156 29764 204212 29766
rect 204260 29818 204316 29820
rect 204260 29766 204262 29818
rect 204262 29766 204314 29818
rect 204314 29766 204316 29818
rect 204260 29764 204316 29766
rect 204364 29818 204420 29820
rect 204364 29766 204366 29818
rect 204366 29766 204418 29818
rect 204418 29766 204420 29818
rect 204364 29764 204420 29766
rect 204156 28250 204212 28252
rect 204156 28198 204158 28250
rect 204158 28198 204210 28250
rect 204210 28198 204212 28250
rect 204156 28196 204212 28198
rect 204260 28250 204316 28252
rect 204260 28198 204262 28250
rect 204262 28198 204314 28250
rect 204314 28198 204316 28250
rect 204260 28196 204316 28198
rect 204364 28250 204420 28252
rect 204364 28198 204366 28250
rect 204366 28198 204418 28250
rect 204418 28198 204420 28250
rect 204364 28196 204420 28198
rect 204156 26682 204212 26684
rect 204156 26630 204158 26682
rect 204158 26630 204210 26682
rect 204210 26630 204212 26682
rect 204156 26628 204212 26630
rect 204260 26682 204316 26684
rect 204260 26630 204262 26682
rect 204262 26630 204314 26682
rect 204314 26630 204316 26682
rect 204260 26628 204316 26630
rect 204364 26682 204420 26684
rect 204364 26630 204366 26682
rect 204366 26630 204418 26682
rect 204418 26630 204420 26682
rect 204364 26628 204420 26630
rect 204156 25114 204212 25116
rect 204156 25062 204158 25114
rect 204158 25062 204210 25114
rect 204210 25062 204212 25114
rect 204156 25060 204212 25062
rect 204260 25114 204316 25116
rect 204260 25062 204262 25114
rect 204262 25062 204314 25114
rect 204314 25062 204316 25114
rect 204260 25060 204316 25062
rect 204364 25114 204420 25116
rect 204364 25062 204366 25114
rect 204366 25062 204418 25114
rect 204418 25062 204420 25114
rect 204364 25060 204420 25062
rect 204156 23546 204212 23548
rect 204156 23494 204158 23546
rect 204158 23494 204210 23546
rect 204210 23494 204212 23546
rect 204156 23492 204212 23494
rect 204260 23546 204316 23548
rect 204260 23494 204262 23546
rect 204262 23494 204314 23546
rect 204314 23494 204316 23546
rect 204260 23492 204316 23494
rect 204364 23546 204420 23548
rect 204364 23494 204366 23546
rect 204366 23494 204418 23546
rect 204418 23494 204420 23546
rect 204364 23492 204420 23494
rect 204156 21978 204212 21980
rect 204156 21926 204158 21978
rect 204158 21926 204210 21978
rect 204210 21926 204212 21978
rect 204156 21924 204212 21926
rect 204260 21978 204316 21980
rect 204260 21926 204262 21978
rect 204262 21926 204314 21978
rect 204314 21926 204316 21978
rect 204260 21924 204316 21926
rect 204364 21978 204420 21980
rect 204364 21926 204366 21978
rect 204366 21926 204418 21978
rect 204418 21926 204420 21978
rect 204364 21924 204420 21926
rect 204156 20410 204212 20412
rect 204156 20358 204158 20410
rect 204158 20358 204210 20410
rect 204210 20358 204212 20410
rect 204156 20356 204212 20358
rect 204260 20410 204316 20412
rect 204260 20358 204262 20410
rect 204262 20358 204314 20410
rect 204314 20358 204316 20410
rect 204260 20356 204316 20358
rect 204364 20410 204420 20412
rect 204364 20358 204366 20410
rect 204366 20358 204418 20410
rect 204418 20358 204420 20410
rect 204364 20356 204420 20358
rect 204156 18842 204212 18844
rect 204156 18790 204158 18842
rect 204158 18790 204210 18842
rect 204210 18790 204212 18842
rect 204156 18788 204212 18790
rect 204260 18842 204316 18844
rect 204260 18790 204262 18842
rect 204262 18790 204314 18842
rect 204314 18790 204316 18842
rect 204260 18788 204316 18790
rect 204364 18842 204420 18844
rect 204364 18790 204366 18842
rect 204366 18790 204418 18842
rect 204418 18790 204420 18842
rect 204364 18788 204420 18790
rect 197260 17612 197316 17668
rect 204156 17274 204212 17276
rect 204156 17222 204158 17274
rect 204158 17222 204210 17274
rect 204210 17222 204212 17274
rect 204156 17220 204212 17222
rect 204260 17274 204316 17276
rect 204260 17222 204262 17274
rect 204262 17222 204314 17274
rect 204314 17222 204316 17274
rect 204260 17220 204316 17222
rect 204364 17274 204420 17276
rect 204364 17222 204366 17274
rect 204366 17222 204418 17274
rect 204418 17222 204420 17274
rect 204364 17220 204420 17222
rect 204156 15706 204212 15708
rect 204156 15654 204158 15706
rect 204158 15654 204210 15706
rect 204210 15654 204212 15706
rect 204156 15652 204212 15654
rect 204260 15706 204316 15708
rect 204260 15654 204262 15706
rect 204262 15654 204314 15706
rect 204314 15654 204316 15706
rect 204260 15652 204316 15654
rect 204364 15706 204420 15708
rect 204364 15654 204366 15706
rect 204366 15654 204418 15706
rect 204418 15654 204420 15706
rect 204364 15652 204420 15654
rect 204156 14138 204212 14140
rect 204156 14086 204158 14138
rect 204158 14086 204210 14138
rect 204210 14086 204212 14138
rect 204156 14084 204212 14086
rect 204260 14138 204316 14140
rect 204260 14086 204262 14138
rect 204262 14086 204314 14138
rect 204314 14086 204316 14138
rect 204260 14084 204316 14086
rect 204364 14138 204420 14140
rect 204364 14086 204366 14138
rect 204366 14086 204418 14138
rect 204418 14086 204420 14138
rect 204364 14084 204420 14086
rect 193116 12796 193172 12852
rect 204156 12570 204212 12572
rect 204156 12518 204158 12570
rect 204158 12518 204210 12570
rect 204210 12518 204212 12570
rect 204156 12516 204212 12518
rect 204260 12570 204316 12572
rect 204260 12518 204262 12570
rect 204262 12518 204314 12570
rect 204314 12518 204316 12570
rect 204260 12516 204316 12518
rect 204364 12570 204420 12572
rect 204364 12518 204366 12570
rect 204366 12518 204418 12570
rect 204418 12518 204420 12570
rect 204364 12516 204420 12518
rect 188796 11786 188852 11788
rect 188796 11734 188798 11786
rect 188798 11734 188850 11786
rect 188850 11734 188852 11786
rect 188796 11732 188852 11734
rect 188900 11786 188956 11788
rect 188900 11734 188902 11786
rect 188902 11734 188954 11786
rect 188954 11734 188956 11786
rect 188900 11732 188956 11734
rect 189004 11786 189060 11788
rect 189004 11734 189006 11786
rect 189006 11734 189058 11786
rect 189058 11734 189060 11786
rect 189004 11732 189060 11734
rect 204156 11002 204212 11004
rect 204156 10950 204158 11002
rect 204158 10950 204210 11002
rect 204210 10950 204212 11002
rect 204156 10948 204212 10950
rect 204260 11002 204316 11004
rect 204260 10950 204262 11002
rect 204262 10950 204314 11002
rect 204314 10950 204316 11002
rect 204260 10948 204316 10950
rect 204364 11002 204420 11004
rect 204364 10950 204366 11002
rect 204366 10950 204418 11002
rect 204418 10950 204420 11002
rect 204364 10948 204420 10950
rect 188796 10218 188852 10220
rect 188796 10166 188798 10218
rect 188798 10166 188850 10218
rect 188850 10166 188852 10218
rect 188796 10164 188852 10166
rect 188900 10218 188956 10220
rect 188900 10166 188902 10218
rect 188902 10166 188954 10218
rect 188954 10166 188956 10218
rect 188900 10164 188956 10166
rect 189004 10218 189060 10220
rect 189004 10166 189006 10218
rect 189006 10166 189058 10218
rect 189058 10166 189060 10218
rect 189004 10164 189060 10166
rect 204156 9434 204212 9436
rect 204156 9382 204158 9434
rect 204158 9382 204210 9434
rect 204210 9382 204212 9434
rect 204156 9380 204212 9382
rect 204260 9434 204316 9436
rect 204260 9382 204262 9434
rect 204262 9382 204314 9434
rect 204314 9382 204316 9434
rect 204260 9380 204316 9382
rect 204364 9434 204420 9436
rect 204364 9382 204366 9434
rect 204366 9382 204418 9434
rect 204418 9382 204420 9434
rect 204364 9380 204420 9382
rect 188796 8650 188852 8652
rect 188796 8598 188798 8650
rect 188798 8598 188850 8650
rect 188850 8598 188852 8650
rect 188796 8596 188852 8598
rect 188900 8650 188956 8652
rect 188900 8598 188902 8650
rect 188902 8598 188954 8650
rect 188954 8598 188956 8650
rect 188900 8596 188956 8598
rect 189004 8650 189060 8652
rect 189004 8598 189006 8650
rect 189006 8598 189058 8650
rect 189058 8598 189060 8650
rect 189004 8596 189060 8598
rect 204156 7866 204212 7868
rect 204156 7814 204158 7866
rect 204158 7814 204210 7866
rect 204210 7814 204212 7866
rect 204156 7812 204212 7814
rect 204260 7866 204316 7868
rect 204260 7814 204262 7866
rect 204262 7814 204314 7866
rect 204314 7814 204316 7866
rect 204260 7812 204316 7814
rect 204364 7866 204420 7868
rect 204364 7814 204366 7866
rect 204366 7814 204418 7866
rect 204418 7814 204420 7866
rect 204364 7812 204420 7814
rect 217532 46002 217588 46004
rect 217532 45950 217534 46002
rect 217534 45950 217586 46002
rect 217586 45950 217588 46002
rect 217532 45948 217588 45950
rect 209356 14252 209412 14308
rect 213948 12684 214004 12740
rect 205772 7644 205828 7700
rect 188796 7082 188852 7084
rect 188796 7030 188798 7082
rect 188798 7030 188850 7082
rect 188850 7030 188852 7082
rect 188796 7028 188852 7030
rect 188900 7082 188956 7084
rect 188900 7030 188902 7082
rect 188902 7030 188954 7082
rect 188954 7030 188956 7082
rect 188900 7028 188956 7030
rect 189004 7082 189060 7084
rect 189004 7030 189006 7082
rect 189006 7030 189058 7082
rect 189058 7030 189060 7082
rect 189004 7028 189060 7030
rect 213948 6860 214004 6916
rect 204156 6298 204212 6300
rect 204156 6246 204158 6298
rect 204158 6246 204210 6298
rect 204210 6246 204212 6298
rect 204156 6244 204212 6246
rect 204260 6298 204316 6300
rect 204260 6246 204262 6298
rect 204262 6246 204314 6298
rect 204314 6246 204316 6298
rect 204260 6244 204316 6246
rect 204364 6298 204420 6300
rect 204364 6246 204366 6298
rect 204366 6246 204418 6298
rect 204418 6246 204420 6298
rect 204364 6244 204420 6246
rect 189308 6076 189364 6132
rect 188796 5514 188852 5516
rect 188796 5462 188798 5514
rect 188798 5462 188850 5514
rect 188850 5462 188852 5514
rect 188796 5460 188852 5462
rect 188900 5514 188956 5516
rect 188900 5462 188902 5514
rect 188902 5462 188954 5514
rect 188954 5462 188956 5514
rect 188900 5460 188956 5462
rect 189004 5514 189060 5516
rect 189004 5462 189006 5514
rect 189006 5462 189058 5514
rect 189058 5462 189060 5514
rect 189004 5460 189060 5462
rect 184492 4172 184548 4228
rect 182252 2380 182308 2436
rect 188796 3946 188852 3948
rect 188796 3894 188798 3946
rect 188798 3894 188850 3946
rect 188850 3894 188852 3946
rect 188796 3892 188852 3894
rect 188900 3946 188956 3948
rect 188900 3894 188902 3946
rect 188902 3894 188954 3946
rect 188954 3894 188956 3946
rect 188900 3892 188956 3894
rect 189004 3946 189060 3948
rect 189004 3894 189006 3946
rect 189006 3894 189058 3946
rect 189058 3894 189060 3946
rect 189004 3892 189060 3894
rect 186620 3724 186676 3780
rect 186396 3442 186452 3444
rect 186396 3390 186398 3442
rect 186398 3390 186450 3442
rect 186450 3390 186452 3442
rect 186396 3388 186452 3390
rect 186844 3388 186900 3444
rect 192108 5964 192164 6020
rect 194684 5628 194740 5684
rect 194460 3442 194516 3444
rect 194460 3390 194462 3442
rect 194462 3390 194514 3442
rect 194514 3390 194516 3442
rect 194460 3388 194516 3390
rect 204156 4730 204212 4732
rect 204156 4678 204158 4730
rect 204158 4678 204210 4730
rect 204210 4678 204212 4730
rect 204156 4676 204212 4678
rect 204260 4730 204316 4732
rect 204260 4678 204262 4730
rect 204262 4678 204314 4730
rect 204314 4678 204316 4730
rect 204260 4676 204316 4678
rect 204364 4730 204420 4732
rect 204364 4678 204366 4730
rect 204366 4678 204418 4730
rect 204418 4678 204420 4730
rect 204364 4676 204420 4678
rect 211596 3666 211652 3668
rect 211596 3614 211598 3666
rect 211598 3614 211650 3666
rect 211650 3614 211652 3666
rect 211596 3612 211652 3614
rect 216636 4508 216692 4564
rect 195020 3442 195076 3444
rect 195020 3390 195022 3442
rect 195022 3390 195074 3442
rect 195074 3390 195076 3442
rect 195020 3388 195076 3390
rect 197932 2156 197988 2212
rect 200620 1372 200676 1428
rect 204156 3162 204212 3164
rect 204156 3110 204158 3162
rect 204158 3110 204210 3162
rect 204210 3110 204212 3162
rect 204156 3108 204212 3110
rect 204260 3162 204316 3164
rect 204260 3110 204262 3162
rect 204262 3110 204314 3162
rect 204314 3110 204316 3162
rect 204260 3108 204316 3110
rect 204364 3162 204420 3164
rect 204364 3110 204366 3162
rect 204366 3110 204418 3162
rect 204418 3110 204420 3162
rect 204364 3108 204420 3110
rect 203980 1596 204036 1652
rect 205996 3276 206052 3332
rect 208684 1484 208740 1540
<< metal3 >>
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 65906 46228 65916 46284
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 66180 46228 66190 46284
rect 96626 46228 96636 46284
rect 96692 46228 96740 46284
rect 96796 46228 96844 46284
rect 96900 46228 96910 46284
rect 127346 46228 127356 46284
rect 127412 46228 127460 46284
rect 127516 46228 127564 46284
rect 127620 46228 127630 46284
rect 158066 46228 158076 46284
rect 158132 46228 158180 46284
rect 158236 46228 158284 46284
rect 158340 46228 158350 46284
rect 188786 46228 188796 46284
rect 188852 46228 188900 46284
rect 188956 46228 189004 46284
rect 189060 46228 189070 46284
rect 148082 46060 148092 46116
rect 148148 46060 150444 46116
rect 150500 46060 150510 46116
rect 31602 45948 31612 46004
rect 31668 45948 32172 46004
rect 32228 45948 32238 46004
rect 150322 45948 150332 46004
rect 150388 45948 205212 46004
rect 205268 45948 205278 46004
rect 205762 45948 205772 46004
rect 205828 45948 217532 46004
rect 217588 45948 217598 46004
rect 19842 45836 19852 45892
rect 19908 45836 22652 45892
rect 22708 45836 22718 45892
rect 36530 45836 36540 45892
rect 36596 45836 37772 45892
rect 37828 45836 37838 45892
rect 44146 45836 44156 45892
rect 44212 45836 47852 45892
rect 47908 45836 47918 45892
rect 54114 45836 54124 45892
rect 54180 45836 55132 45892
rect 55188 45836 58044 45892
rect 58100 45836 58110 45892
rect 100146 45836 100156 45892
rect 100212 45836 100828 45892
rect 100884 45836 100894 45892
rect 103954 45836 103964 45892
rect 104020 45836 104636 45892
rect 104692 45836 104702 45892
rect 172498 45836 172508 45892
rect 172564 45836 173292 45892
rect 173348 45836 173358 45892
rect 176306 45836 176316 45892
rect 176372 45836 177100 45892
rect 177156 45836 177166 45892
rect 184034 45836 184044 45892
rect 184100 45836 184828 45892
rect 184884 45836 184894 45892
rect 65874 45724 65884 45780
rect 65940 45724 66556 45780
rect 66612 45724 130172 45780
rect 130228 45724 130238 45780
rect 187282 45724 187292 45780
rect 187348 45724 189196 45780
rect 189252 45724 189262 45780
rect 196532 45724 201292 45780
rect 201348 45724 201358 45780
rect 50082 45612 50092 45668
rect 50148 45612 50540 45668
rect 50596 45612 52892 45668
rect 52948 45612 52958 45668
rect 58146 45612 58156 45668
rect 58212 45612 58940 45668
rect 58996 45612 61292 45668
rect 61348 45612 61358 45668
rect 62066 45612 62076 45668
rect 62132 45612 62748 45668
rect 62804 45612 69692 45668
rect 69748 45612 69758 45668
rect 69906 45612 69916 45668
rect 69972 45612 70364 45668
rect 70420 45612 73276 45668
rect 73332 45612 73342 45668
rect 73490 45612 73500 45668
rect 73556 45612 74172 45668
rect 74228 45612 76412 45668
rect 76468 45612 76478 45668
rect 139906 45612 139916 45668
rect 139972 45612 144284 45668
rect 144340 45612 144350 45668
rect 196532 45556 196588 45724
rect 182242 45500 182252 45556
rect 182308 45500 196588 45556
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 50546 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50830 45500
rect 81266 45444 81276 45500
rect 81332 45444 81380 45500
rect 81436 45444 81484 45500
rect 81540 45444 81550 45500
rect 111986 45444 111996 45500
rect 112052 45444 112100 45500
rect 112156 45444 112204 45500
rect 112260 45444 112270 45500
rect 142706 45444 142716 45500
rect 142772 45444 142820 45500
rect 142876 45444 142924 45500
rect 142980 45444 142990 45500
rect 173426 45444 173436 45500
rect 173492 45444 173540 45500
rect 173596 45444 173644 45500
rect 173700 45444 173710 45500
rect 204146 45444 204156 45500
rect 204212 45444 204260 45500
rect 204316 45444 204364 45500
rect 204420 45444 204430 45500
rect 32722 45388 32732 45444
rect 32788 45388 42812 45444
rect 42868 45388 42878 45444
rect 152114 45276 152124 45332
rect 152180 45276 153356 45332
rect 153412 45276 153422 45332
rect 135650 45164 135660 45220
rect 135716 45164 140588 45220
rect 140644 45164 140654 45220
rect 12338 45052 12348 45108
rect 12404 45052 126028 45108
rect 125972 44996 126028 45052
rect 125972 44940 138124 44996
rect 138180 44940 139804 44996
rect 139860 44940 139870 44996
rect 141922 44940 141932 44996
rect 141988 44940 152124 44996
rect 152180 44940 152190 44996
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 65906 44660 65916 44716
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 66180 44660 66190 44716
rect 96626 44660 96636 44716
rect 96692 44660 96740 44716
rect 96796 44660 96844 44716
rect 96900 44660 96910 44716
rect 127346 44660 127356 44716
rect 127412 44660 127460 44716
rect 127516 44660 127564 44716
rect 127620 44660 127630 44716
rect 158066 44660 158076 44716
rect 158132 44660 158180 44716
rect 158236 44660 158284 44716
rect 158340 44660 158350 44716
rect 188786 44660 188796 44716
rect 188852 44660 188900 44716
rect 188956 44660 189004 44716
rect 189060 44660 189070 44716
rect 131954 44268 131964 44324
rect 132020 44268 135100 44324
rect 135156 44268 135166 44324
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 50546 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50830 43932
rect 81266 43876 81276 43932
rect 81332 43876 81380 43932
rect 81436 43876 81484 43932
rect 81540 43876 81550 43932
rect 111986 43876 111996 43932
rect 112052 43876 112100 43932
rect 112156 43876 112204 43932
rect 112260 43876 112270 43932
rect 142706 43876 142716 43932
rect 142772 43876 142820 43932
rect 142876 43876 142924 43932
rect 142980 43876 142990 43932
rect 173426 43876 173436 43932
rect 173492 43876 173540 43932
rect 173596 43876 173644 43932
rect 173700 43876 173710 43932
rect 204146 43876 204156 43932
rect 204212 43876 204260 43932
rect 204316 43876 204364 43932
rect 204420 43876 204430 43932
rect 167122 43708 167132 43764
rect 167188 43708 173068 43764
rect 173124 43708 173134 43764
rect 80098 43596 80108 43652
rect 80164 43596 126028 43652
rect 125972 43540 126028 43596
rect 125972 43484 135772 43540
rect 135828 43484 136108 43540
rect 136164 43484 136174 43540
rect 137228 43484 138684 43540
rect 138740 43484 140364 43540
rect 140420 43484 140430 43540
rect 137228 43428 137284 43484
rect 135090 43372 135100 43428
rect 135156 43372 135996 43428
rect 136052 43372 137228 43428
rect 137284 43372 137294 43428
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 65906 43092 65916 43148
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 66180 43092 66190 43148
rect 96626 43092 96636 43148
rect 96692 43092 96740 43148
rect 96796 43092 96844 43148
rect 96900 43092 96910 43148
rect 127346 43092 127356 43148
rect 127412 43092 127460 43148
rect 127516 43092 127564 43148
rect 127620 43092 127630 43148
rect 158066 43092 158076 43148
rect 158132 43092 158180 43148
rect 158236 43092 158284 43148
rect 158340 43092 158350 43148
rect 188786 43092 188796 43148
rect 188852 43092 188900 43148
rect 188956 43092 189004 43148
rect 189060 43092 189070 43148
rect 137554 42924 137564 42980
rect 137620 42924 138124 42980
rect 138180 42924 138190 42980
rect 134754 42700 134764 42756
rect 134820 42700 137900 42756
rect 137956 42700 137966 42756
rect 136210 42476 136220 42532
rect 136276 42476 137788 42532
rect 137844 42476 137854 42532
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 50546 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50830 42364
rect 81266 42308 81276 42364
rect 81332 42308 81380 42364
rect 81436 42308 81484 42364
rect 81540 42308 81550 42364
rect 111986 42308 111996 42364
rect 112052 42308 112100 42364
rect 112156 42308 112204 42364
rect 112260 42308 112270 42364
rect 142706 42308 142716 42364
rect 142772 42308 142820 42364
rect 142876 42308 142924 42364
rect 142980 42308 142990 42364
rect 173426 42308 173436 42364
rect 173492 42308 173540 42364
rect 173596 42308 173644 42364
rect 173700 42308 173710 42364
rect 204146 42308 204156 42364
rect 204212 42308 204260 42364
rect 204316 42308 204364 42364
rect 204420 42308 204430 42364
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 65906 41524 65916 41580
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 66180 41524 66190 41580
rect 96626 41524 96636 41580
rect 96692 41524 96740 41580
rect 96796 41524 96844 41580
rect 96900 41524 96910 41580
rect 127346 41524 127356 41580
rect 127412 41524 127460 41580
rect 127516 41524 127564 41580
rect 127620 41524 127630 41580
rect 158066 41524 158076 41580
rect 158132 41524 158180 41580
rect 158236 41524 158284 41580
rect 158340 41524 158350 41580
rect 188786 41524 188796 41580
rect 188852 41524 188900 41580
rect 188956 41524 189004 41580
rect 189060 41524 189070 41580
rect 92194 41132 92204 41188
rect 92260 41132 118412 41188
rect 118468 41132 118478 41188
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 50546 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50830 40796
rect 81266 40740 81276 40796
rect 81332 40740 81380 40796
rect 81436 40740 81484 40796
rect 81540 40740 81550 40796
rect 111986 40740 111996 40796
rect 112052 40740 112100 40796
rect 112156 40740 112204 40796
rect 112260 40740 112270 40796
rect 142706 40740 142716 40796
rect 142772 40740 142820 40796
rect 142876 40740 142924 40796
rect 142980 40740 142990 40796
rect 173426 40740 173436 40796
rect 173492 40740 173540 40796
rect 173596 40740 173644 40796
rect 173700 40740 173710 40796
rect 204146 40740 204156 40796
rect 204212 40740 204260 40796
rect 204316 40740 204364 40796
rect 204420 40740 204430 40796
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 65906 39956 65916 40012
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 66180 39956 66190 40012
rect 96626 39956 96636 40012
rect 96692 39956 96740 40012
rect 96796 39956 96844 40012
rect 96900 39956 96910 40012
rect 127346 39956 127356 40012
rect 127412 39956 127460 40012
rect 127516 39956 127564 40012
rect 127620 39956 127630 40012
rect 158066 39956 158076 40012
rect 158132 39956 158180 40012
rect 158236 39956 158284 40012
rect 158340 39956 158350 40012
rect 188786 39956 188796 40012
rect 188852 39956 188900 40012
rect 188956 39956 189004 40012
rect 189060 39956 189070 40012
rect 88162 39452 88172 39508
rect 88228 39452 133980 39508
rect 134036 39452 134046 39508
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 50546 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50830 39228
rect 81266 39172 81276 39228
rect 81332 39172 81380 39228
rect 81436 39172 81484 39228
rect 81540 39172 81550 39228
rect 111986 39172 111996 39228
rect 112052 39172 112100 39228
rect 112156 39172 112204 39228
rect 112260 39172 112270 39228
rect 142706 39172 142716 39228
rect 142772 39172 142820 39228
rect 142876 39172 142924 39228
rect 142980 39172 142990 39228
rect 173426 39172 173436 39228
rect 173492 39172 173540 39228
rect 173596 39172 173644 39228
rect 173700 39172 173710 39228
rect 204146 39172 204156 39228
rect 204212 39172 204260 39228
rect 204316 39172 204364 39228
rect 204420 39172 204430 39228
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 65906 38388 65916 38444
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 66180 38388 66190 38444
rect 96626 38388 96636 38444
rect 96692 38388 96740 38444
rect 96796 38388 96844 38444
rect 96900 38388 96910 38444
rect 127346 38388 127356 38444
rect 127412 38388 127460 38444
rect 127516 38388 127564 38444
rect 127620 38388 127630 38444
rect 158066 38388 158076 38444
rect 158132 38388 158180 38444
rect 158236 38388 158284 38444
rect 158340 38388 158350 38444
rect 188786 38388 188796 38444
rect 188852 38388 188900 38444
rect 188956 38388 189004 38444
rect 189060 38388 189070 38444
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 50546 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50830 37660
rect 81266 37604 81276 37660
rect 81332 37604 81380 37660
rect 81436 37604 81484 37660
rect 81540 37604 81550 37660
rect 111986 37604 111996 37660
rect 112052 37604 112100 37660
rect 112156 37604 112204 37660
rect 112260 37604 112270 37660
rect 142706 37604 142716 37660
rect 142772 37604 142820 37660
rect 142876 37604 142924 37660
rect 142980 37604 142990 37660
rect 173426 37604 173436 37660
rect 173492 37604 173540 37660
rect 173596 37604 173644 37660
rect 173700 37604 173710 37660
rect 204146 37604 204156 37660
rect 204212 37604 204260 37660
rect 204316 37604 204364 37660
rect 204420 37604 204430 37660
rect 2930 37100 2940 37156
rect 2996 37100 118748 37156
rect 118804 37100 119308 37156
rect 119364 37100 119374 37156
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 65906 36820 65916 36876
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 66180 36820 66190 36876
rect 96626 36820 96636 36876
rect 96692 36820 96740 36876
rect 96796 36820 96844 36876
rect 96900 36820 96910 36876
rect 127346 36820 127356 36876
rect 127412 36820 127460 36876
rect 127516 36820 127564 36876
rect 127620 36820 127630 36876
rect 158066 36820 158076 36876
rect 158132 36820 158180 36876
rect 158236 36820 158284 36876
rect 158340 36820 158350 36876
rect 188786 36820 188796 36876
rect 188852 36820 188900 36876
rect 188956 36820 189004 36876
rect 189060 36820 189070 36876
rect 117170 36204 117180 36260
rect 117236 36204 124236 36260
rect 124292 36204 130508 36260
rect 130564 36204 131068 36260
rect 131124 36204 131134 36260
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 50546 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50830 36092
rect 81266 36036 81276 36092
rect 81332 36036 81380 36092
rect 81436 36036 81484 36092
rect 81540 36036 81550 36092
rect 111986 36036 111996 36092
rect 112052 36036 112100 36092
rect 112156 36036 112204 36092
rect 112260 36036 112270 36092
rect 142706 36036 142716 36092
rect 142772 36036 142820 36092
rect 142876 36036 142924 36092
rect 142980 36036 142990 36092
rect 173426 36036 173436 36092
rect 173492 36036 173540 36092
rect 173596 36036 173644 36092
rect 173700 36036 173710 36092
rect 204146 36036 204156 36092
rect 204212 36036 204260 36092
rect 204316 36036 204364 36092
rect 204420 36036 204430 36092
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 65906 35252 65916 35308
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 66180 35252 66190 35308
rect 96626 35252 96636 35308
rect 96692 35252 96740 35308
rect 96796 35252 96844 35308
rect 96900 35252 96910 35308
rect 127346 35252 127356 35308
rect 127412 35252 127460 35308
rect 127516 35252 127564 35308
rect 127620 35252 127630 35308
rect 158066 35252 158076 35308
rect 158132 35252 158180 35308
rect 158236 35252 158284 35308
rect 158340 35252 158350 35308
rect 188786 35252 188796 35308
rect 188852 35252 188900 35308
rect 188956 35252 189004 35308
rect 189060 35252 189070 35308
rect 136098 35196 136108 35252
rect 136164 35196 136780 35252
rect 136836 35196 136846 35252
rect 84130 34636 84140 34692
rect 84196 34636 132636 34692
rect 132692 34636 132702 34692
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 50546 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50830 34524
rect 81266 34468 81276 34524
rect 81332 34468 81380 34524
rect 81436 34468 81484 34524
rect 81540 34468 81550 34524
rect 111986 34468 111996 34524
rect 112052 34468 112100 34524
rect 112156 34468 112204 34524
rect 112260 34468 112270 34524
rect 142706 34468 142716 34524
rect 142772 34468 142820 34524
rect 142876 34468 142924 34524
rect 142980 34468 142990 34524
rect 173426 34468 173436 34524
rect 173492 34468 173540 34524
rect 173596 34468 173644 34524
rect 173700 34468 173710 34524
rect 204146 34468 204156 34524
rect 204212 34468 204260 34524
rect 204316 34468 204364 34524
rect 204420 34468 204430 34524
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 65906 33684 65916 33740
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 66180 33684 66190 33740
rect 96626 33684 96636 33740
rect 96692 33684 96740 33740
rect 96796 33684 96844 33740
rect 96900 33684 96910 33740
rect 127346 33684 127356 33740
rect 127412 33684 127460 33740
rect 127516 33684 127564 33740
rect 127620 33684 127630 33740
rect 158066 33684 158076 33740
rect 158132 33684 158180 33740
rect 158236 33684 158284 33740
rect 158340 33684 158350 33740
rect 188786 33684 188796 33740
rect 188852 33684 188900 33740
rect 188956 33684 189004 33740
rect 189060 33684 189070 33740
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 50546 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50830 32956
rect 81266 32900 81276 32956
rect 81332 32900 81380 32956
rect 81436 32900 81484 32956
rect 81540 32900 81550 32956
rect 111986 32900 111996 32956
rect 112052 32900 112100 32956
rect 112156 32900 112204 32956
rect 112260 32900 112270 32956
rect 142706 32900 142716 32956
rect 142772 32900 142820 32956
rect 142876 32900 142924 32956
rect 142980 32900 142990 32956
rect 173426 32900 173436 32956
rect 173492 32900 173540 32956
rect 173596 32900 173644 32956
rect 173700 32900 173710 32956
rect 204146 32900 204156 32956
rect 204212 32900 204260 32956
rect 204316 32900 204364 32956
rect 204420 32900 204430 32956
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 65906 32116 65916 32172
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 66180 32116 66190 32172
rect 96626 32116 96636 32172
rect 96692 32116 96740 32172
rect 96796 32116 96844 32172
rect 96900 32116 96910 32172
rect 127346 32116 127356 32172
rect 127412 32116 127460 32172
rect 127516 32116 127564 32172
rect 127620 32116 127630 32172
rect 158066 32116 158076 32172
rect 158132 32116 158180 32172
rect 158236 32116 158284 32172
rect 158340 32116 158350 32172
rect 188786 32116 188796 32172
rect 188852 32116 188900 32172
rect 188956 32116 189004 32172
rect 189060 32116 189070 32172
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 50546 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50830 31388
rect 81266 31332 81276 31388
rect 81332 31332 81380 31388
rect 81436 31332 81484 31388
rect 81540 31332 81550 31388
rect 111986 31332 111996 31388
rect 112052 31332 112100 31388
rect 112156 31332 112204 31388
rect 112260 31332 112270 31388
rect 142706 31332 142716 31388
rect 142772 31332 142820 31388
rect 142876 31332 142924 31388
rect 142980 31332 142990 31388
rect 173426 31332 173436 31388
rect 173492 31332 173540 31388
rect 173596 31332 173644 31388
rect 173700 31332 173710 31388
rect 204146 31332 204156 31388
rect 204212 31332 204260 31388
rect 204316 31332 204364 31388
rect 204420 31332 204430 31388
rect 106530 30828 106540 30884
rect 106596 30828 108220 30884
rect 108276 30828 109900 30884
rect 109956 30828 109966 30884
rect 113586 30828 113596 30884
rect 113652 30828 116732 30884
rect 116788 30828 117628 30884
rect 117684 30828 117694 30884
rect 118402 30828 118412 30884
rect 118468 30828 136332 30884
rect 136388 30828 138124 30884
rect 138180 30828 138190 30884
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 65906 30548 65916 30604
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 66180 30548 66190 30604
rect 96626 30548 96636 30604
rect 96692 30548 96740 30604
rect 96796 30548 96844 30604
rect 96900 30548 96910 30604
rect 127346 30548 127356 30604
rect 127412 30548 127460 30604
rect 127516 30548 127564 30604
rect 127620 30548 127630 30604
rect 158066 30548 158076 30604
rect 158132 30548 158180 30604
rect 158236 30548 158284 30604
rect 158340 30548 158350 30604
rect 188786 30548 188796 30604
rect 188852 30548 188900 30604
rect 188956 30548 189004 30604
rect 189060 30548 189070 30604
rect 104972 30268 108892 30324
rect 108948 30268 113372 30324
rect 113428 30268 113438 30324
rect 104972 30212 105028 30268
rect 112364 30212 112420 30268
rect 96226 30156 96236 30212
rect 96292 30156 96684 30212
rect 96740 30156 101276 30212
rect 101332 30156 104412 30212
rect 104468 30156 104972 30212
rect 105028 30156 105038 30212
rect 112354 30156 112364 30212
rect 112420 30156 112430 30212
rect 125346 30156 125356 30212
rect 125412 30156 128940 30212
rect 128996 30156 129948 30212
rect 130004 30156 132860 30212
rect 132916 30156 134428 30212
rect 134484 30156 136220 30212
rect 136276 30156 136780 30212
rect 136836 30156 136846 30212
rect 93762 30044 93772 30100
rect 93828 30044 95452 30100
rect 95508 30044 97132 30100
rect 97188 30044 97198 30100
rect 101602 30044 101612 30100
rect 101668 30044 103740 30100
rect 103796 30044 105420 30100
rect 105476 30044 105486 30100
rect 110786 30044 110796 30100
rect 110852 30044 111692 30100
rect 111748 30044 112924 30100
rect 112980 30044 112990 30100
rect 126130 30044 126140 30100
rect 126196 30044 128268 30100
rect 128324 30044 129500 30100
rect 129556 30044 129566 30100
rect 132626 30044 132636 30100
rect 132692 30044 133644 30100
rect 133700 30044 133710 30100
rect 118738 29932 118748 29988
rect 118804 29932 120428 29988
rect 120484 29932 121324 29988
rect 121380 29932 121390 29988
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 50546 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50830 29820
rect 81266 29764 81276 29820
rect 81332 29764 81380 29820
rect 81436 29764 81484 29820
rect 81540 29764 81550 29820
rect 111986 29764 111996 29820
rect 112052 29764 112100 29820
rect 112156 29764 112204 29820
rect 112260 29764 112270 29820
rect 142706 29764 142716 29820
rect 142772 29764 142820 29820
rect 142876 29764 142924 29820
rect 142980 29764 142990 29820
rect 173426 29764 173436 29820
rect 173492 29764 173540 29820
rect 173596 29764 173644 29820
rect 173700 29764 173710 29820
rect 204146 29764 204156 29820
rect 204212 29764 204260 29820
rect 204316 29764 204364 29820
rect 204420 29764 204430 29820
rect 124450 29596 124460 29652
rect 124516 29596 125356 29652
rect 125412 29596 125422 29652
rect 133970 29596 133980 29652
rect 134036 29596 135772 29652
rect 135828 29596 135838 29652
rect 97906 29260 97916 29316
rect 97972 29260 100044 29316
rect 100100 29260 101724 29316
rect 101780 29260 101790 29316
rect 121762 29260 121772 29316
rect 121828 29260 123676 29316
rect 123732 29260 124908 29316
rect 124964 29260 124974 29316
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 65906 28980 65916 29036
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 66180 28980 66190 29036
rect 96626 28980 96636 29036
rect 96692 28980 96740 29036
rect 96796 28980 96844 29036
rect 96900 28980 96910 29036
rect 127346 28980 127356 29036
rect 127412 28980 127460 29036
rect 127516 28980 127564 29036
rect 127620 28980 127630 29036
rect 158066 28980 158076 29036
rect 158132 28980 158180 29036
rect 158236 28980 158284 29036
rect 158340 28980 158350 29036
rect 188786 28980 188796 29036
rect 188852 28980 188900 29036
rect 188956 28980 189004 29036
rect 189060 28980 189070 29036
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 50546 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50830 28252
rect 81266 28196 81276 28252
rect 81332 28196 81380 28252
rect 81436 28196 81484 28252
rect 81540 28196 81550 28252
rect 111986 28196 111996 28252
rect 112052 28196 112100 28252
rect 112156 28196 112204 28252
rect 112260 28196 112270 28252
rect 142706 28196 142716 28252
rect 142772 28196 142820 28252
rect 142876 28196 142924 28252
rect 142980 28196 142990 28252
rect 173426 28196 173436 28252
rect 173492 28196 173540 28252
rect 173596 28196 173644 28252
rect 173700 28196 173710 28252
rect 204146 28196 204156 28252
rect 204212 28196 204260 28252
rect 204316 28196 204364 28252
rect 204420 28196 204430 28252
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 65906 27412 65916 27468
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 66180 27412 66190 27468
rect 96626 27412 96636 27468
rect 96692 27412 96740 27468
rect 96796 27412 96844 27468
rect 96900 27412 96910 27468
rect 127346 27412 127356 27468
rect 127412 27412 127460 27468
rect 127516 27412 127564 27468
rect 127620 27412 127630 27468
rect 158066 27412 158076 27468
rect 158132 27412 158180 27468
rect 158236 27412 158284 27468
rect 158340 27412 158350 27468
rect 188786 27412 188796 27468
rect 188852 27412 188900 27468
rect 188956 27412 189004 27468
rect 189060 27412 189070 27468
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 50546 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50830 26684
rect 81266 26628 81276 26684
rect 81332 26628 81380 26684
rect 81436 26628 81484 26684
rect 81540 26628 81550 26684
rect 111986 26628 111996 26684
rect 112052 26628 112100 26684
rect 112156 26628 112204 26684
rect 112260 26628 112270 26684
rect 142706 26628 142716 26684
rect 142772 26628 142820 26684
rect 142876 26628 142924 26684
rect 142980 26628 142990 26684
rect 173426 26628 173436 26684
rect 173492 26628 173540 26684
rect 173596 26628 173644 26684
rect 173700 26628 173710 26684
rect 204146 26628 204156 26684
rect 204212 26628 204260 26684
rect 204316 26628 204364 26684
rect 204420 26628 204430 26684
rect 23874 26012 23884 26068
rect 23940 26012 55132 26068
rect 55188 26012 55198 26068
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 65906 25844 65916 25900
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 66180 25844 66190 25900
rect 96626 25844 96636 25900
rect 96692 25844 96740 25900
rect 96796 25844 96844 25900
rect 96900 25844 96910 25900
rect 127346 25844 127356 25900
rect 127412 25844 127460 25900
rect 127516 25844 127564 25900
rect 127620 25844 127630 25900
rect 158066 25844 158076 25900
rect 158132 25844 158180 25900
rect 158236 25844 158284 25900
rect 158340 25844 158350 25900
rect 188786 25844 188796 25900
rect 188852 25844 188900 25900
rect 188956 25844 189004 25900
rect 189060 25844 189070 25900
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 50546 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50830 25116
rect 81266 25060 81276 25116
rect 81332 25060 81380 25116
rect 81436 25060 81484 25116
rect 81540 25060 81550 25116
rect 111986 25060 111996 25116
rect 112052 25060 112100 25116
rect 112156 25060 112204 25116
rect 112260 25060 112270 25116
rect 142706 25060 142716 25116
rect 142772 25060 142820 25116
rect 142876 25060 142924 25116
rect 142980 25060 142990 25116
rect 173426 25060 173436 25116
rect 173492 25060 173540 25116
rect 173596 25060 173644 25116
rect 173700 25060 173710 25116
rect 204146 25060 204156 25116
rect 204212 25060 204260 25116
rect 204316 25060 204364 25116
rect 204420 25060 204430 25116
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 65906 24276 65916 24332
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 66180 24276 66190 24332
rect 96626 24276 96636 24332
rect 96692 24276 96740 24332
rect 96796 24276 96844 24332
rect 96900 24276 96910 24332
rect 127346 24276 127356 24332
rect 127412 24276 127460 24332
rect 127516 24276 127564 24332
rect 127620 24276 127630 24332
rect 158066 24276 158076 24332
rect 158132 24276 158180 24332
rect 158236 24276 158284 24332
rect 158340 24276 158350 24332
rect 188786 24276 188796 24332
rect 188852 24276 188900 24332
rect 188956 24276 189004 24332
rect 189060 24276 189070 24332
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 50546 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50830 23548
rect 81266 23492 81276 23548
rect 81332 23492 81380 23548
rect 81436 23492 81484 23548
rect 81540 23492 81550 23548
rect 111986 23492 111996 23548
rect 112052 23492 112100 23548
rect 112156 23492 112204 23548
rect 112260 23492 112270 23548
rect 142706 23492 142716 23548
rect 142772 23492 142820 23548
rect 142876 23492 142924 23548
rect 142980 23492 142990 23548
rect 173426 23492 173436 23548
rect 173492 23492 173540 23548
rect 173596 23492 173644 23548
rect 173700 23492 173710 23548
rect 204146 23492 204156 23548
rect 204212 23492 204260 23548
rect 204316 23492 204364 23548
rect 204420 23492 204430 23548
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 65906 22708 65916 22764
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 66180 22708 66190 22764
rect 96626 22708 96636 22764
rect 96692 22708 96740 22764
rect 96796 22708 96844 22764
rect 96900 22708 96910 22764
rect 127346 22708 127356 22764
rect 127412 22708 127460 22764
rect 127516 22708 127564 22764
rect 127620 22708 127630 22764
rect 158066 22708 158076 22764
rect 158132 22708 158180 22764
rect 158236 22708 158284 22764
rect 158340 22708 158350 22764
rect 188786 22708 188796 22764
rect 188852 22708 188900 22764
rect 188956 22708 189004 22764
rect 189060 22708 189070 22764
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 50546 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50830 21980
rect 81266 21924 81276 21980
rect 81332 21924 81380 21980
rect 81436 21924 81484 21980
rect 81540 21924 81550 21980
rect 111986 21924 111996 21980
rect 112052 21924 112100 21980
rect 112156 21924 112204 21980
rect 112260 21924 112270 21980
rect 142706 21924 142716 21980
rect 142772 21924 142820 21980
rect 142876 21924 142924 21980
rect 142980 21924 142990 21980
rect 173426 21924 173436 21980
rect 173492 21924 173540 21980
rect 173596 21924 173644 21980
rect 173700 21924 173710 21980
rect 204146 21924 204156 21980
rect 204212 21924 204260 21980
rect 204316 21924 204364 21980
rect 204420 21924 204430 21980
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 65906 21140 65916 21196
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 66180 21140 66190 21196
rect 96626 21140 96636 21196
rect 96692 21140 96740 21196
rect 96796 21140 96844 21196
rect 96900 21140 96910 21196
rect 127346 21140 127356 21196
rect 127412 21140 127460 21196
rect 127516 21140 127564 21196
rect 127620 21140 127630 21196
rect 158066 21140 158076 21196
rect 158132 21140 158180 21196
rect 158236 21140 158284 21196
rect 158340 21140 158350 21196
rect 188786 21140 188796 21196
rect 188852 21140 188900 21196
rect 188956 21140 189004 21196
rect 189060 21140 189070 21196
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 50546 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50830 20412
rect 81266 20356 81276 20412
rect 81332 20356 81380 20412
rect 81436 20356 81484 20412
rect 81540 20356 81550 20412
rect 111986 20356 111996 20412
rect 112052 20356 112100 20412
rect 112156 20356 112204 20412
rect 112260 20356 112270 20412
rect 142706 20356 142716 20412
rect 142772 20356 142820 20412
rect 142876 20356 142924 20412
rect 142980 20356 142990 20412
rect 173426 20356 173436 20412
rect 173492 20356 173540 20412
rect 173596 20356 173644 20412
rect 173700 20356 173710 20412
rect 204146 20356 204156 20412
rect 204212 20356 204260 20412
rect 204316 20356 204364 20412
rect 204420 20356 204430 20412
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 65906 19572 65916 19628
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 66180 19572 66190 19628
rect 96626 19572 96636 19628
rect 96692 19572 96740 19628
rect 96796 19572 96844 19628
rect 96900 19572 96910 19628
rect 127346 19572 127356 19628
rect 127412 19572 127460 19628
rect 127516 19572 127564 19628
rect 127620 19572 127630 19628
rect 158066 19572 158076 19628
rect 158132 19572 158180 19628
rect 158236 19572 158284 19628
rect 158340 19572 158350 19628
rect 188786 19572 188796 19628
rect 188852 19572 188900 19628
rect 188956 19572 189004 19628
rect 189060 19572 189070 19628
rect 47842 19292 47852 19348
rect 47908 19292 68572 19348
rect 68628 19292 68638 19348
rect 76402 19292 76412 19348
rect 76468 19292 136220 19348
rect 136276 19292 136286 19348
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 50546 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50830 18844
rect 81266 18788 81276 18844
rect 81332 18788 81380 18844
rect 81436 18788 81484 18844
rect 81540 18788 81550 18844
rect 111986 18788 111996 18844
rect 112052 18788 112100 18844
rect 112156 18788 112204 18844
rect 112260 18788 112270 18844
rect 142706 18788 142716 18844
rect 142772 18788 142820 18844
rect 142876 18788 142924 18844
rect 142980 18788 142990 18844
rect 173426 18788 173436 18844
rect 173492 18788 173540 18844
rect 173596 18788 173644 18844
rect 173700 18788 173710 18844
rect 204146 18788 204156 18844
rect 204212 18788 204260 18844
rect 204316 18788 204364 18844
rect 204420 18788 204430 18844
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 65906 18004 65916 18060
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 66180 18004 66190 18060
rect 96626 18004 96636 18060
rect 96692 18004 96740 18060
rect 96796 18004 96844 18060
rect 96900 18004 96910 18060
rect 127346 18004 127356 18060
rect 127412 18004 127460 18060
rect 127516 18004 127564 18060
rect 127620 18004 127630 18060
rect 158066 18004 158076 18060
rect 158132 18004 158180 18060
rect 158236 18004 158284 18060
rect 158340 18004 158350 18060
rect 188786 18004 188796 18060
rect 188852 18004 188900 18060
rect 188956 18004 189004 18060
rect 189060 18004 189070 18060
rect 73266 17612 73276 17668
rect 73332 17612 134652 17668
rect 134708 17612 134718 17668
rect 145842 17612 145852 17668
rect 145908 17612 197260 17668
rect 197316 17612 197326 17668
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 50546 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50830 17276
rect 81266 17220 81276 17276
rect 81332 17220 81380 17276
rect 81436 17220 81484 17276
rect 81540 17220 81550 17276
rect 111986 17220 111996 17276
rect 112052 17220 112100 17276
rect 112156 17220 112204 17276
rect 112260 17220 112270 17276
rect 142706 17220 142716 17276
rect 142772 17220 142820 17276
rect 142876 17220 142924 17276
rect 142980 17220 142990 17276
rect 173426 17220 173436 17276
rect 173492 17220 173540 17276
rect 173596 17220 173644 17276
rect 173700 17220 173710 17276
rect 204146 17220 204156 17276
rect 204212 17220 204260 17276
rect 204316 17220 204364 17276
rect 204420 17220 204430 17276
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 65906 16436 65916 16492
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 66180 16436 66190 16492
rect 96626 16436 96636 16492
rect 96692 16436 96740 16492
rect 96796 16436 96844 16492
rect 96900 16436 96910 16492
rect 127346 16436 127356 16492
rect 127412 16436 127460 16492
rect 127516 16436 127564 16492
rect 127620 16436 127630 16492
rect 158066 16436 158076 16492
rect 158132 16436 158180 16492
rect 158236 16436 158284 16492
rect 158340 16436 158350 16492
rect 188786 16436 188796 16492
rect 188852 16436 188900 16492
rect 188956 16436 189004 16492
rect 189060 16436 189070 16492
rect 37762 15932 37772 15988
rect 37828 15932 63196 15988
rect 63252 15932 63262 15988
rect 69682 15932 69692 15988
rect 69748 15932 132748 15988
rect 132804 15932 132814 15988
rect 162866 15932 162876 15988
rect 162932 15932 184604 15988
rect 184660 15932 184670 15988
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 50546 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50830 15708
rect 81266 15652 81276 15708
rect 81332 15652 81380 15708
rect 81436 15652 81484 15708
rect 81540 15652 81550 15708
rect 111986 15652 111996 15708
rect 112052 15652 112100 15708
rect 112156 15652 112204 15708
rect 112260 15652 112270 15708
rect 142706 15652 142716 15708
rect 142772 15652 142820 15708
rect 142876 15652 142924 15708
rect 142980 15652 142990 15708
rect 173426 15652 173436 15708
rect 173492 15652 173540 15708
rect 173596 15652 173644 15708
rect 173700 15652 173710 15708
rect 204146 15652 204156 15708
rect 204212 15652 204260 15708
rect 204316 15652 204364 15708
rect 204420 15652 204430 15708
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 65906 14868 65916 14924
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 66180 14868 66190 14924
rect 96626 14868 96636 14924
rect 96692 14868 96740 14924
rect 96796 14868 96844 14924
rect 96900 14868 96910 14924
rect 127346 14868 127356 14924
rect 127412 14868 127460 14924
rect 127516 14868 127564 14924
rect 127620 14868 127630 14924
rect 158066 14868 158076 14924
rect 158132 14868 158180 14924
rect 158236 14868 158284 14924
rect 158340 14868 158350 14924
rect 188786 14868 188796 14924
rect 188852 14868 188900 14924
rect 188956 14868 189004 14924
rect 189060 14868 189070 14924
rect 168018 14364 168028 14420
rect 168084 14364 180684 14420
rect 180740 14364 180750 14420
rect 42802 14252 42812 14308
rect 42868 14252 59948 14308
rect 60004 14252 60014 14308
rect 61282 14252 61292 14308
rect 61348 14252 138012 14308
rect 138068 14252 138078 14308
rect 153682 14252 153692 14308
rect 153748 14252 209356 14308
rect 209412 14252 209422 14308
rect 164658 14140 164668 14196
rect 164724 14140 169260 14196
rect 169316 14140 169326 14196
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 50546 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50830 14140
rect 81266 14084 81276 14140
rect 81332 14084 81380 14140
rect 81436 14084 81484 14140
rect 81540 14084 81550 14140
rect 111986 14084 111996 14140
rect 112052 14084 112100 14140
rect 112156 14084 112204 14140
rect 112260 14084 112270 14140
rect 142706 14084 142716 14140
rect 142772 14084 142820 14140
rect 142876 14084 142924 14140
rect 142980 14084 142990 14140
rect 173426 14084 173436 14140
rect 173492 14084 173540 14140
rect 173596 14084 173644 14140
rect 173700 14084 173710 14140
rect 204146 14084 204156 14140
rect 204212 14084 204260 14140
rect 204316 14084 204364 14140
rect 204420 14084 204430 14140
rect 140242 13468 140252 13524
rect 140308 13468 148204 13524
rect 148260 13468 148270 13524
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 65906 13300 65916 13356
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 66180 13300 66190 13356
rect 96626 13300 96636 13356
rect 96692 13300 96740 13356
rect 96796 13300 96844 13356
rect 96900 13300 96910 13356
rect 127346 13300 127356 13356
rect 127412 13300 127460 13356
rect 127516 13300 127564 13356
rect 127620 13300 127630 13356
rect 158066 13300 158076 13356
rect 158132 13300 158180 13356
rect 158236 13300 158284 13356
rect 158340 13300 158350 13356
rect 188786 13300 188796 13356
rect 188852 13300 188900 13356
rect 188956 13300 189004 13356
rect 189060 13300 189070 13356
rect 143602 12908 143612 12964
rect 143668 12908 187292 12964
rect 187348 12908 187358 12964
rect 146402 12796 146412 12852
rect 146468 12796 193116 12852
rect 193172 12796 193182 12852
rect 28914 12684 28924 12740
rect 28980 12684 57820 12740
rect 57876 12684 57886 12740
rect 58034 12684 58044 12740
rect 58100 12684 140140 12740
rect 140196 12684 140206 12740
rect 153234 12684 153244 12740
rect 153300 12684 154588 12740
rect 154644 12684 154654 12740
rect 156212 12684 213948 12740
rect 214004 12684 214014 12740
rect 156212 12628 156268 12684
rect 150770 12572 150780 12628
rect 150836 12572 156268 12628
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 50546 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50830 12572
rect 81266 12516 81276 12572
rect 81332 12516 81380 12572
rect 81436 12516 81484 12572
rect 81540 12516 81550 12572
rect 111986 12516 111996 12572
rect 112052 12516 112100 12572
rect 112156 12516 112204 12572
rect 112260 12516 112270 12572
rect 142706 12516 142716 12572
rect 142772 12516 142820 12572
rect 142876 12516 142924 12572
rect 142980 12516 142990 12572
rect 173426 12516 173436 12572
rect 173492 12516 173540 12572
rect 173596 12516 173644 12572
rect 173700 12516 173710 12572
rect 204146 12516 204156 12572
rect 204212 12516 204260 12572
rect 204316 12516 204364 12572
rect 204420 12516 204430 12572
rect 163314 12012 163324 12068
rect 163380 12012 176876 12068
rect 176932 12012 176942 12068
rect 159852 11788 164444 11844
rect 164500 11788 164510 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 65906 11732 65916 11788
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 66180 11732 66190 11788
rect 96626 11732 96636 11788
rect 96692 11732 96740 11788
rect 96796 11732 96844 11788
rect 96900 11732 96910 11788
rect 127346 11732 127356 11788
rect 127412 11732 127460 11788
rect 127516 11732 127564 11788
rect 127620 11732 127630 11788
rect 158066 11732 158076 11788
rect 158132 11732 158180 11788
rect 158236 11732 158284 11788
rect 158340 11732 158350 11788
rect 147746 11676 147756 11732
rect 147812 11676 150332 11732
rect 150388 11676 150398 11732
rect 159852 11620 159908 11788
rect 188786 11732 188796 11788
rect 188852 11732 188900 11788
rect 188956 11732 189004 11788
rect 189060 11732 189070 11788
rect 160738 11676 160748 11732
rect 160804 11676 162876 11732
rect 162932 11676 162942 11732
rect 167972 11620 168028 11732
rect 168084 11676 168094 11732
rect 139122 11564 139132 11620
rect 139188 11564 150500 11620
rect 157154 11564 157164 11620
rect 157220 11564 157724 11620
rect 157780 11564 159908 11620
rect 162978 11564 162988 11620
rect 163044 11564 168028 11620
rect 137890 11452 137900 11508
rect 137956 11452 146860 11508
rect 146916 11452 147308 11508
rect 147364 11452 149212 11508
rect 149268 11452 149278 11508
rect 150444 11284 150500 11564
rect 150658 11452 150668 11508
rect 150724 11452 156492 11508
rect 156548 11452 160300 11508
rect 160356 11452 160366 11508
rect 156034 11340 156044 11396
rect 156100 11340 156716 11396
rect 156772 11340 156782 11396
rect 163986 11340 163996 11396
rect 164052 11340 164668 11396
rect 164724 11340 164734 11396
rect 40226 11228 40236 11284
rect 40292 11228 65436 11284
rect 65492 11228 65502 11284
rect 77858 11228 77868 11284
rect 77924 11228 131068 11284
rect 131124 11228 131134 11284
rect 150444 11228 156268 11284
rect 156212 11172 156268 11228
rect 52882 11116 52892 11172
rect 52948 11116 140028 11172
rect 140084 11116 140094 11172
rect 156212 11116 159852 11172
rect 159908 11116 159918 11172
rect 162642 11116 162652 11172
rect 162708 11116 163548 11172
rect 163604 11116 163614 11172
rect 144452 11004 156716 11060
rect 156772 11004 156782 11060
rect 156940 11004 162876 11060
rect 162932 11004 163772 11060
rect 163828 11004 163838 11060
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 50546 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50830 11004
rect 81266 10948 81276 11004
rect 81332 10948 81380 11004
rect 81436 10948 81484 11004
rect 81540 10948 81550 11004
rect 111986 10948 111996 11004
rect 112052 10948 112100 11004
rect 112156 10948 112204 11004
rect 112260 10948 112270 11004
rect 142706 10948 142716 11004
rect 142772 10948 142820 11004
rect 142876 10948 142924 11004
rect 142980 10948 142990 11004
rect 144452 10836 144508 11004
rect 156940 10948 156996 11004
rect 173426 10948 173436 11004
rect 173492 10948 173540 11004
rect 173596 10948 173644 11004
rect 173700 10948 173710 11004
rect 204146 10948 204156 11004
rect 204212 10948 204260 11004
rect 204316 10948 204364 11004
rect 204420 10948 204430 11004
rect 155138 10892 155148 10948
rect 155204 10892 156940 10948
rect 156996 10892 157006 10948
rect 161970 10892 161980 10948
rect 162036 10892 162988 10948
rect 163044 10892 163054 10948
rect 138450 10780 138460 10836
rect 138516 10780 144508 10836
rect 147858 10780 147868 10836
rect 147924 10780 148204 10836
rect 148260 10780 148270 10836
rect 161522 10780 161532 10836
rect 161588 10780 162316 10836
rect 162372 10780 162382 10836
rect 163986 10780 163996 10836
rect 164052 10780 164444 10836
rect 164500 10780 167132 10836
rect 167188 10780 167198 10836
rect 154018 10668 154028 10724
rect 154084 10668 154924 10724
rect 154980 10668 154990 10724
rect 156212 10668 160524 10724
rect 160580 10668 162092 10724
rect 162148 10668 162158 10724
rect 149650 10556 149660 10612
rect 149716 10556 151228 10612
rect 151284 10556 151294 10612
rect 156212 10500 156268 10668
rect 160290 10556 160300 10612
rect 160356 10556 161196 10612
rect 161252 10556 161262 10612
rect 162530 10556 162540 10612
rect 162596 10556 163324 10612
rect 163380 10556 163390 10612
rect 135874 10444 135884 10500
rect 135940 10444 146188 10500
rect 146244 10444 147532 10500
rect 147588 10444 148204 10500
rect 148260 10444 148270 10500
rect 153570 10444 153580 10500
rect 153636 10444 155596 10500
rect 155652 10444 156268 10500
rect 156706 10444 156716 10500
rect 156772 10444 161644 10500
rect 161700 10444 161710 10500
rect 137666 10332 137676 10388
rect 137732 10332 152236 10388
rect 152292 10332 152302 10388
rect 148866 10220 148876 10276
rect 148932 10220 150556 10276
rect 150612 10220 153132 10276
rect 153188 10220 154812 10276
rect 154868 10220 154878 10276
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 65906 10164 65916 10220
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 66180 10164 66190 10220
rect 96626 10164 96636 10220
rect 96692 10164 96740 10220
rect 96796 10164 96844 10220
rect 96900 10164 96910 10220
rect 127346 10164 127356 10220
rect 127412 10164 127460 10220
rect 127516 10164 127564 10220
rect 127620 10164 127630 10220
rect 158066 10164 158076 10220
rect 158132 10164 158180 10220
rect 158236 10164 158284 10220
rect 158340 10164 158350 10220
rect 188786 10164 188796 10220
rect 188852 10164 188900 10220
rect 188956 10164 189004 10220
rect 189060 10164 189070 10220
rect 138226 10108 138236 10164
rect 138292 10108 139132 10164
rect 139188 10108 139198 10164
rect 139356 10108 151452 10164
rect 151508 10108 151518 10164
rect 158508 10108 160412 10164
rect 160468 10108 160478 10164
rect 139356 10052 139412 10108
rect 158508 10052 158564 10108
rect 138674 9996 138684 10052
rect 138740 9996 139412 10052
rect 155586 9996 155596 10052
rect 155652 9996 157164 10052
rect 157220 9996 158564 10052
rect 112578 9884 112588 9940
rect 112644 9884 153244 9940
rect 153300 9884 153310 9940
rect 148754 9772 148764 9828
rect 148820 9772 149548 9828
rect 149604 9772 150108 9828
rect 150164 9772 151564 9828
rect 151620 9772 151630 9828
rect 156034 9772 156044 9828
rect 156100 9772 156110 9828
rect 156258 9772 156268 9828
rect 156324 9772 156828 9828
rect 156884 9772 156894 9828
rect 156044 9716 156100 9772
rect 114482 9660 114492 9716
rect 114548 9660 151732 9716
rect 156044 9660 157052 9716
rect 157108 9660 157118 9716
rect 151676 9604 151732 9660
rect 147970 9548 147980 9604
rect 148036 9548 148652 9604
rect 148708 9548 150668 9604
rect 150724 9548 150734 9604
rect 151666 9548 151676 9604
rect 151732 9548 151742 9604
rect 155698 9548 155708 9604
rect 155764 9548 157276 9604
rect 157332 9548 157342 9604
rect 146066 9436 146076 9492
rect 146132 9436 150108 9492
rect 150164 9436 150780 9492
rect 150836 9436 150846 9492
rect 156044 9436 160076 9492
rect 160132 9436 161532 9492
rect 161588 9436 161598 9492
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 50546 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50830 9436
rect 81266 9380 81276 9436
rect 81332 9380 81380 9436
rect 81436 9380 81484 9436
rect 81540 9380 81550 9436
rect 111986 9380 111996 9436
rect 112052 9380 112100 9436
rect 112156 9380 112204 9436
rect 112260 9380 112270 9436
rect 142706 9380 142716 9436
rect 142772 9380 142820 9436
rect 142876 9380 142924 9436
rect 142980 9380 142990 9436
rect 156044 9268 156100 9436
rect 173426 9380 173436 9436
rect 173492 9380 173540 9436
rect 173596 9380 173644 9436
rect 173700 9380 173710 9436
rect 204146 9380 204156 9436
rect 204212 9380 204260 9436
rect 204316 9380 204364 9436
rect 204420 9380 204430 9436
rect 22642 9212 22652 9268
rect 22708 9212 52108 9268
rect 52164 9212 52174 9268
rect 140914 9212 140924 9268
rect 140980 9212 141932 9268
rect 141988 9212 141998 9268
rect 148418 9212 148428 9268
rect 148484 9212 149772 9268
rect 149828 9212 151116 9268
rect 151172 9212 151182 9268
rect 152114 9212 152124 9268
rect 152180 9212 156044 9268
rect 156100 9212 156110 9268
rect 131058 9100 131068 9156
rect 131124 9100 135324 9156
rect 135380 9100 135390 9156
rect 135986 9100 135996 9156
rect 136052 9100 138124 9156
rect 138180 9100 138684 9156
rect 138740 9100 138750 9156
rect 139122 9100 139132 9156
rect 139188 9100 139804 9156
rect 139860 9100 140252 9156
rect 140308 9100 140318 9156
rect 148530 9100 148540 9156
rect 148596 9100 149324 9156
rect 149380 9100 149390 9156
rect 110338 8988 110348 9044
rect 110404 8988 134540 9044
rect 134596 8988 135548 9044
rect 135604 8988 135614 9044
rect 152450 8988 152460 9044
rect 152516 8988 153916 9044
rect 153972 8988 153982 9044
rect 149650 8876 149660 8932
rect 149716 8876 160636 8932
rect 160692 8876 160702 8932
rect 153458 8764 153468 8820
rect 153524 8764 156828 8820
rect 156884 8764 156894 8820
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 65906 8596 65916 8652
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 66180 8596 66190 8652
rect 96626 8596 96636 8652
rect 96692 8596 96740 8652
rect 96796 8596 96844 8652
rect 96900 8596 96910 8652
rect 127346 8596 127356 8652
rect 127412 8596 127460 8652
rect 127516 8596 127564 8652
rect 127620 8596 127630 8652
rect 158066 8596 158076 8652
rect 158132 8596 158180 8652
rect 158236 8596 158284 8652
rect 158340 8596 158350 8652
rect 188786 8596 188796 8652
rect 188852 8596 188900 8652
rect 188956 8596 189004 8652
rect 189060 8596 189070 8652
rect 144452 8540 155428 8596
rect 162754 8540 162764 8596
rect 162820 8540 163996 8596
rect 164052 8540 164062 8596
rect 144452 8484 144508 8540
rect 155372 8484 155428 8540
rect 88050 8428 88060 8484
rect 88116 8428 144508 8484
rect 151666 8428 151676 8484
rect 151732 8428 152796 8484
rect 152852 8428 152862 8484
rect 153234 8428 153244 8484
rect 153300 8428 153804 8484
rect 153860 8428 153870 8484
rect 155362 8428 155372 8484
rect 155428 8428 155438 8484
rect 161186 8428 161196 8484
rect 161252 8428 163436 8484
rect 163492 8428 163502 8484
rect 130162 8316 130172 8372
rect 130228 8316 132860 8372
rect 132916 8316 132926 8372
rect 147858 8316 147868 8372
rect 147924 8316 148540 8372
rect 148596 8316 156828 8372
rect 156884 8316 156894 8372
rect 134306 8204 134316 8260
rect 134372 8204 139468 8260
rect 139524 8204 139534 8260
rect 150994 8204 151004 8260
rect 151060 8204 152348 8260
rect 152404 8204 159292 8260
rect 159348 8204 162428 8260
rect 162484 8204 162494 8260
rect 135762 8092 135772 8148
rect 135828 8092 136332 8148
rect 136388 8092 136398 8148
rect 142146 8092 142156 8148
rect 142212 8092 156380 8148
rect 156436 8092 156446 8148
rect 135538 7980 135548 8036
rect 135604 7980 145292 8036
rect 145348 7980 145358 8036
rect 162754 7980 162764 8036
rect 162820 7980 164332 8036
rect 164388 7980 164398 8036
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 50546 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50830 7868
rect 81266 7812 81276 7868
rect 81332 7812 81380 7868
rect 81436 7812 81484 7868
rect 81540 7812 81550 7868
rect 111986 7812 111996 7868
rect 112052 7812 112100 7868
rect 112156 7812 112204 7868
rect 112260 7812 112270 7868
rect 142706 7812 142716 7868
rect 142772 7812 142820 7868
rect 142876 7812 142924 7868
rect 142980 7812 142990 7868
rect 173426 7812 173436 7868
rect 173492 7812 173540 7868
rect 173596 7812 173644 7868
rect 173700 7812 173710 7868
rect 204146 7812 204156 7868
rect 204212 7812 204260 7868
rect 204316 7812 204364 7868
rect 204420 7812 204430 7868
rect 151890 7756 151900 7812
rect 151956 7756 153132 7812
rect 153188 7756 160076 7812
rect 160132 7756 160142 7812
rect 140802 7644 140812 7700
rect 140868 7644 142940 7700
rect 142996 7644 143006 7700
rect 143266 7644 143276 7700
rect 143332 7644 145740 7700
rect 145796 7644 145806 7700
rect 147858 7644 147868 7700
rect 147924 7644 147934 7700
rect 155138 7644 155148 7700
rect 155204 7644 205772 7700
rect 205828 7644 205838 7700
rect 147868 7588 147924 7644
rect 15810 7532 15820 7588
rect 15876 7532 49756 7588
rect 49812 7532 49822 7588
rect 132514 7532 132524 7588
rect 132580 7532 133196 7588
rect 133252 7532 134540 7588
rect 134596 7532 135660 7588
rect 135716 7532 135726 7588
rect 137666 7532 137676 7588
rect 137732 7532 147924 7588
rect 161746 7532 161756 7588
rect 161812 7532 162204 7588
rect 162260 7532 162988 7588
rect 163044 7532 163054 7588
rect 130498 7420 130508 7476
rect 130564 7420 131740 7476
rect 131796 7420 131806 7476
rect 131954 7420 131964 7476
rect 132020 7420 135548 7476
rect 135604 7420 135614 7476
rect 139234 7420 139244 7476
rect 139300 7420 140588 7476
rect 140644 7420 140654 7476
rect 144050 7420 144060 7476
rect 144116 7420 148204 7476
rect 148260 7420 148270 7476
rect 148754 7420 148764 7476
rect 148820 7420 150892 7476
rect 150948 7420 151228 7476
rect 151284 7420 151294 7476
rect 152114 7420 152124 7476
rect 152180 7420 152908 7476
rect 152964 7420 153580 7476
rect 153636 7420 153646 7476
rect 162530 7420 162540 7476
rect 162596 7420 168028 7476
rect 167972 7364 168028 7420
rect 148866 7308 148876 7364
rect 148932 7308 151116 7364
rect 151172 7308 152236 7364
rect 152292 7308 152302 7364
rect 152450 7308 152460 7364
rect 152516 7308 154924 7364
rect 154980 7308 154990 7364
rect 160290 7308 160300 7364
rect 160356 7308 161084 7364
rect 161140 7308 161420 7364
rect 161476 7308 161486 7364
rect 167972 7308 170492 7364
rect 170548 7308 170558 7364
rect 149986 7196 149996 7252
rect 150052 7196 155148 7252
rect 155204 7196 155214 7252
rect 156594 7196 156604 7252
rect 156660 7196 161644 7252
rect 161700 7196 161710 7252
rect 145170 7084 145180 7140
rect 145236 7084 145404 7140
rect 145460 7084 150220 7140
rect 150276 7084 152124 7140
rect 152180 7084 152190 7140
rect 162428 7084 162652 7140
rect 162708 7084 162718 7140
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 65906 7028 65916 7084
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 66180 7028 66190 7084
rect 96626 7028 96636 7084
rect 96692 7028 96740 7084
rect 96796 7028 96844 7084
rect 96900 7028 96910 7084
rect 127346 7028 127356 7084
rect 127412 7028 127460 7084
rect 127516 7028 127564 7084
rect 127620 7028 127630 7084
rect 158066 7028 158076 7084
rect 158132 7028 158180 7084
rect 158236 7028 158284 7084
rect 158340 7028 158350 7084
rect 162428 7028 162484 7084
rect 188786 7028 188796 7084
rect 188852 7028 188900 7084
rect 188956 7028 189004 7084
rect 189060 7028 189070 7084
rect 147634 6972 147644 7028
rect 147700 6972 150108 7028
rect 150164 6972 156268 7028
rect 162418 6972 162428 7028
rect 162484 6972 162494 7028
rect 162726 6972 162764 7028
rect 162820 6972 162830 7028
rect 156212 6916 156268 6972
rect 33170 6860 33180 6916
rect 33236 6860 97468 6916
rect 97524 6860 97534 6916
rect 131730 6860 131740 6916
rect 131796 6860 133084 6916
rect 133140 6860 133150 6916
rect 134194 6860 134204 6916
rect 134260 6860 145180 6916
rect 145236 6860 145246 6916
rect 151442 6860 151452 6916
rect 151508 6860 151518 6916
rect 154242 6860 154252 6916
rect 154308 6860 155820 6916
rect 155876 6860 155886 6916
rect 156212 6860 213948 6916
rect 214004 6860 214014 6916
rect 151452 6804 151508 6860
rect 39218 6748 39228 6804
rect 39284 6748 105532 6804
rect 105588 6748 105598 6804
rect 137218 6748 137228 6804
rect 137284 6748 139468 6804
rect 139524 6748 139534 6804
rect 145058 6748 145068 6804
rect 145124 6748 148092 6804
rect 148148 6748 148158 6804
rect 151452 6748 156268 6804
rect 160514 6748 160524 6804
rect 160580 6748 161532 6804
rect 161588 6748 161598 6804
rect 163314 6748 163324 6804
rect 163380 6748 167804 6804
rect 167860 6748 167870 6804
rect 156212 6692 156268 6748
rect 131282 6636 131292 6692
rect 131348 6636 133084 6692
rect 133140 6636 133150 6692
rect 135538 6636 135548 6692
rect 135604 6636 136332 6692
rect 136388 6636 138236 6692
rect 138292 6636 138302 6692
rect 142482 6636 142492 6692
rect 142548 6636 145852 6692
rect 145908 6636 145918 6692
rect 151106 6636 151116 6692
rect 151172 6636 154700 6692
rect 154756 6636 154766 6692
rect 156212 6636 159628 6692
rect 159684 6636 159694 6692
rect 160962 6636 160972 6692
rect 161028 6636 161196 6692
rect 161252 6636 161262 6692
rect 162642 6636 162652 6692
rect 162708 6636 164220 6692
rect 164276 6636 164286 6692
rect 106754 6524 106764 6580
rect 106820 6524 132076 6580
rect 132132 6524 132142 6580
rect 140354 6524 140364 6580
rect 140420 6524 144620 6580
rect 144676 6524 144686 6580
rect 160066 6524 160076 6580
rect 160132 6524 161420 6580
rect 161476 6524 162876 6580
rect 162932 6524 162942 6580
rect 163090 6524 163100 6580
rect 163156 6524 163884 6580
rect 163940 6524 163950 6580
rect 73042 6412 73052 6468
rect 73108 6412 125580 6468
rect 125636 6412 125646 6468
rect 135762 6412 135772 6468
rect 135828 6412 137900 6468
rect 137956 6412 139356 6468
rect 139412 6412 139422 6468
rect 141810 6412 141820 6468
rect 141876 6412 144284 6468
rect 144340 6412 144350 6468
rect 148978 6412 148988 6468
rect 149044 6412 153244 6468
rect 153300 6412 156044 6468
rect 156100 6412 156110 6468
rect 159618 6412 159628 6468
rect 159684 6412 160748 6468
rect 160804 6412 160814 6468
rect 161634 6412 161644 6468
rect 161700 6412 163772 6468
rect 163828 6412 163838 6468
rect 163986 6412 163996 6468
rect 164052 6412 164090 6468
rect 164546 6412 164556 6468
rect 164612 6412 165116 6468
rect 165172 6412 184828 6468
rect 152674 6300 152684 6356
rect 152740 6300 161980 6356
rect 162036 6300 162046 6356
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 50546 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50830 6300
rect 81266 6244 81276 6300
rect 81332 6244 81380 6300
rect 81436 6244 81484 6300
rect 81540 6244 81550 6300
rect 111986 6244 111996 6300
rect 112052 6244 112100 6300
rect 112156 6244 112204 6300
rect 112260 6244 112270 6300
rect 142706 6244 142716 6300
rect 142772 6244 142820 6300
rect 142876 6244 142924 6300
rect 142980 6244 142990 6300
rect 173426 6244 173436 6300
rect 173492 6244 173540 6300
rect 173596 6244 173644 6300
rect 173700 6244 173710 6300
rect 149650 6188 149660 6244
rect 149716 6188 151452 6244
rect 151508 6188 151518 6244
rect 152562 6188 152572 6244
rect 152628 6188 163324 6244
rect 163380 6188 163390 6244
rect 184772 6132 184828 6412
rect 204146 6244 204156 6300
rect 204212 6244 204260 6300
rect 204316 6244 204364 6300
rect 204420 6244 204430 6300
rect 98578 6076 98588 6132
rect 98644 6076 130060 6132
rect 130116 6076 130126 6132
rect 133746 6076 133756 6132
rect 133812 6076 139132 6132
rect 139188 6076 139198 6132
rect 144452 6076 152460 6132
rect 152516 6076 154028 6132
rect 154084 6076 154094 6132
rect 156818 6076 156828 6132
rect 156884 6076 157948 6132
rect 158004 6076 159964 6132
rect 160020 6076 160300 6132
rect 160356 6076 160366 6132
rect 160738 6076 160748 6132
rect 160804 6076 162764 6132
rect 162820 6076 162830 6132
rect 163510 6076 163548 6132
rect 163604 6076 163614 6132
rect 164210 6076 164220 6132
rect 164276 6076 173068 6132
rect 184772 6076 189308 6132
rect 189364 6076 189374 6132
rect 144452 6020 144508 6076
rect 162764 6020 162820 6076
rect 173012 6020 173068 6076
rect 44482 5964 44492 6020
rect 44548 5964 113372 6020
rect 113428 5964 113438 6020
rect 125122 5964 125132 6020
rect 125188 5964 144508 6020
rect 149874 5964 149884 6020
rect 149940 5964 152124 6020
rect 152180 5964 152190 6020
rect 154802 5964 154812 6020
rect 154868 5964 157724 6020
rect 157780 5964 157790 6020
rect 162764 5964 163996 6020
rect 164052 5964 164062 6020
rect 173012 5964 192108 6020
rect 192164 5964 192174 6020
rect 57026 5852 57036 5908
rect 57092 5852 121212 5908
rect 121268 5852 121278 5908
rect 133970 5852 133980 5908
rect 134036 5852 135100 5908
rect 135156 5852 135166 5908
rect 139122 5852 139132 5908
rect 139188 5852 140644 5908
rect 147298 5852 147308 5908
rect 147364 5852 149436 5908
rect 149492 5852 149502 5908
rect 150098 5852 150108 5908
rect 150164 5852 150668 5908
rect 150724 5852 151340 5908
rect 151396 5852 151900 5908
rect 151956 5852 151966 5908
rect 153682 5852 153692 5908
rect 153748 5852 164108 5908
rect 164164 5852 164174 5908
rect 165106 5852 165116 5908
rect 165172 5852 165564 5908
rect 165620 5852 181244 5908
rect 181300 5852 181310 5908
rect 140588 5796 140644 5852
rect 31490 5740 31500 5796
rect 31556 5740 92764 5796
rect 92820 5740 92830 5796
rect 125972 5740 139468 5796
rect 139524 5740 139534 5796
rect 140578 5740 140588 5796
rect 140644 5740 141036 5796
rect 141092 5740 141102 5796
rect 146066 5740 146076 5796
rect 146132 5740 149100 5796
rect 149156 5740 149166 5796
rect 150210 5740 150220 5796
rect 150276 5740 161868 5796
rect 161924 5740 161934 5796
rect 163762 5740 163772 5796
rect 163828 5740 168028 5796
rect 125972 5684 126028 5740
rect 167972 5684 168028 5740
rect 84242 5628 84252 5684
rect 84308 5628 126028 5684
rect 141810 5628 141820 5684
rect 141876 5628 144284 5684
rect 144340 5628 150332 5684
rect 150388 5628 150398 5684
rect 157154 5628 157164 5684
rect 157220 5628 165004 5684
rect 165060 5628 165070 5684
rect 167972 5628 194684 5684
rect 194740 5628 194750 5684
rect 145730 5516 145740 5572
rect 145796 5516 148540 5572
rect 148596 5516 150556 5572
rect 150612 5516 150622 5572
rect 159730 5516 159740 5572
rect 159796 5516 160748 5572
rect 160804 5516 160814 5572
rect 163762 5516 163772 5572
rect 163828 5516 164556 5572
rect 164612 5516 164622 5572
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 65906 5460 65916 5516
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 66180 5460 66190 5516
rect 96626 5460 96636 5516
rect 96692 5460 96740 5516
rect 96796 5460 96844 5516
rect 96900 5460 96910 5516
rect 127346 5460 127356 5516
rect 127412 5460 127460 5516
rect 127516 5460 127564 5516
rect 127620 5460 127630 5516
rect 158066 5460 158076 5516
rect 158132 5460 158180 5516
rect 158236 5460 158284 5516
rect 158340 5460 158350 5516
rect 188786 5460 188796 5516
rect 188852 5460 188900 5516
rect 188956 5460 189004 5516
rect 189060 5460 189070 5516
rect 141810 5404 141820 5460
rect 141876 5404 145404 5460
rect 145460 5404 145470 5460
rect 153906 5404 153916 5460
rect 153972 5404 154924 5460
rect 154980 5404 155932 5460
rect 155988 5404 155998 5460
rect 161746 5404 161756 5460
rect 161812 5404 162316 5460
rect 162372 5404 163548 5460
rect 163604 5404 164444 5460
rect 164500 5404 164510 5460
rect 89058 5292 89068 5348
rect 89124 5292 133700 5348
rect 135762 5292 135772 5348
rect 135828 5292 136444 5348
rect 136500 5292 136510 5348
rect 141922 5292 141932 5348
rect 141988 5292 153020 5348
rect 153076 5292 153086 5348
rect 155810 5292 155820 5348
rect 155876 5292 156828 5348
rect 156884 5292 156894 5348
rect 157052 5292 157388 5348
rect 157444 5292 157836 5348
rect 157892 5292 157902 5348
rect 159068 5292 162876 5348
rect 162932 5292 162942 5348
rect 163090 5292 163100 5348
rect 163156 5292 164780 5348
rect 164836 5292 165676 5348
rect 165732 5292 165742 5348
rect 133644 5236 133700 5292
rect 157052 5236 157108 5292
rect 5954 5180 5964 5236
rect 6020 5180 6412 5236
rect 6468 5180 7196 5236
rect 7252 5180 7262 5236
rect 59938 5180 59948 5236
rect 60004 5180 60844 5236
rect 60900 5180 60910 5236
rect 93986 5180 93996 5236
rect 94052 5180 109228 5236
rect 109284 5180 109294 5236
rect 109890 5180 109900 5236
rect 109956 5180 110796 5236
rect 110852 5180 110862 5236
rect 113922 5180 113932 5236
rect 113988 5180 114380 5236
rect 114436 5180 116060 5236
rect 116116 5180 116126 5236
rect 116834 5180 116844 5236
rect 116900 5180 133420 5236
rect 133476 5180 133486 5236
rect 133644 5180 137452 5236
rect 137508 5180 137518 5236
rect 142482 5180 142492 5236
rect 142548 5180 145852 5236
rect 145908 5180 145918 5236
rect 152786 5180 152796 5236
rect 152852 5180 153916 5236
rect 153972 5180 153982 5236
rect 156212 5180 157108 5236
rect 157266 5180 157276 5236
rect 157332 5180 157948 5236
rect 158004 5180 158014 5236
rect 156212 5124 156268 5180
rect 159068 5124 159124 5292
rect 161970 5180 161980 5236
rect 162036 5180 163324 5236
rect 163380 5180 163390 5236
rect 163958 5180 163996 5236
rect 164052 5180 164062 5236
rect 165218 5180 165228 5236
rect 165284 5180 166124 5236
rect 166180 5180 166190 5236
rect 108994 5068 109004 5124
rect 109060 5068 110012 5124
rect 110068 5068 110078 5124
rect 138114 5068 138124 5124
rect 138180 5068 140476 5124
rect 140532 5068 141260 5124
rect 141316 5068 141326 5124
rect 142258 5068 142268 5124
rect 142324 5068 143052 5124
rect 143108 5068 143118 5124
rect 144946 5068 144956 5124
rect 145012 5068 146636 5124
rect 146692 5068 148540 5124
rect 148596 5068 148606 5124
rect 154690 5068 154700 5124
rect 154756 5068 155820 5124
rect 155876 5068 156268 5124
rect 156818 5068 156828 5124
rect 156884 5068 159124 5124
rect 159282 5068 159292 5124
rect 159348 5068 160524 5124
rect 160580 5068 160590 5124
rect 161522 5068 161532 5124
rect 161588 5068 166236 5124
rect 166292 5068 166302 5124
rect 135874 4956 135884 5012
rect 135940 4956 138908 5012
rect 138964 4956 138974 5012
rect 141474 4956 141484 5012
rect 141540 4956 147420 5012
rect 147476 4956 147486 5012
rect 151218 4956 151228 5012
rect 151284 4956 152460 5012
rect 152516 4956 156268 5012
rect 156324 4956 156334 5012
rect 156594 4956 156604 5012
rect 156660 4956 158284 5012
rect 158340 4956 161476 5012
rect 162978 4956 162988 5012
rect 163044 4956 178556 5012
rect 178612 4956 178622 5012
rect 161420 4900 161476 4956
rect 46946 4844 46956 4900
rect 47012 4844 117628 4900
rect 117684 4844 117694 4900
rect 136994 4844 137004 4900
rect 137060 4844 138012 4900
rect 138068 4844 138078 4900
rect 138786 4844 138796 4900
rect 138852 4844 140364 4900
rect 140420 4844 140430 4900
rect 142492 4844 146860 4900
rect 146916 4844 146926 4900
rect 150322 4844 150332 4900
rect 150388 4844 153244 4900
rect 153300 4844 153310 4900
rect 154802 4844 154812 4900
rect 154868 4844 157836 4900
rect 157892 4844 157902 4900
rect 158050 4844 158060 4900
rect 158116 4844 159740 4900
rect 159796 4844 159806 4900
rect 161410 4844 161420 4900
rect 161476 4844 163548 4900
rect 163604 4844 163772 4900
rect 163828 4844 163838 4900
rect 142492 4788 142548 4844
rect 135314 4732 135324 4788
rect 135380 4732 142548 4788
rect 144452 4732 150780 4788
rect 150836 4732 150846 4788
rect 157714 4732 157724 4788
rect 157780 4732 168028 4788
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 50546 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50830 4732
rect 81266 4676 81276 4732
rect 81332 4676 81380 4732
rect 81436 4676 81484 4732
rect 81540 4676 81550 4732
rect 111986 4676 111996 4732
rect 112052 4676 112100 4732
rect 112156 4676 112204 4732
rect 112260 4676 112270 4732
rect 142706 4676 142716 4732
rect 142772 4676 142820 4732
rect 142876 4676 142924 4732
rect 142980 4676 142990 4732
rect 144452 4676 144508 4732
rect 127810 4620 127820 4676
rect 127876 4620 137788 4676
rect 137844 4620 137854 4676
rect 138114 4620 138124 4676
rect 138180 4620 139804 4676
rect 139860 4620 139870 4676
rect 143388 4620 144508 4676
rect 149996 4620 152572 4676
rect 152628 4620 155036 4676
rect 155092 4620 155102 4676
rect 161970 4620 161980 4676
rect 162036 4620 164220 4676
rect 164276 4620 164286 4676
rect 143388 4564 143444 4620
rect 35634 4508 35644 4564
rect 35700 4508 101052 4564
rect 101108 4508 101118 4564
rect 130498 4508 130508 4564
rect 130564 4508 143444 4564
rect 149090 4508 149100 4564
rect 149156 4508 149772 4564
rect 149828 4508 149838 4564
rect 149996 4452 150052 4620
rect 167972 4564 168028 4732
rect 173426 4676 173436 4732
rect 173492 4676 173540 4732
rect 173596 4676 173644 4732
rect 173700 4676 173710 4732
rect 204146 4676 204156 4732
rect 204212 4676 204260 4732
rect 204316 4676 204364 4732
rect 204420 4676 204430 4732
rect 153906 4508 153916 4564
rect 153972 4508 155260 4564
rect 155316 4508 155326 4564
rect 161746 4508 161756 4564
rect 161812 4508 163660 4564
rect 163716 4508 163726 4564
rect 167972 4508 216636 4564
rect 216692 4508 216702 4564
rect 51986 4396 51996 4452
rect 52052 4396 52556 4452
rect 52612 4396 73052 4452
rect 73108 4396 73118 4452
rect 77186 4396 77196 4452
rect 77252 4396 136444 4452
rect 136500 4396 136510 4452
rect 137778 4396 137788 4452
rect 137844 4396 150052 4452
rect 150210 4396 150220 4452
rect 150276 4396 162204 4452
rect 162260 4396 162270 4452
rect 162754 4396 162764 4452
rect 162820 4396 165340 4452
rect 165396 4396 165406 4452
rect 55794 4284 55804 4340
rect 55860 4284 57596 4340
rect 57652 4284 57662 4340
rect 66546 4284 66556 4340
rect 66612 4284 68348 4340
rect 68404 4284 68414 4340
rect 78866 4284 78876 4340
rect 78932 4284 79548 4340
rect 79604 4284 80556 4340
rect 80612 4284 80622 4340
rect 81330 4284 81340 4340
rect 81396 4284 84252 4340
rect 84308 4284 84318 4340
rect 87042 4284 87052 4340
rect 87108 4284 88060 4340
rect 88116 4284 88126 4340
rect 93426 4284 93436 4340
rect 93492 4284 132972 4340
rect 133028 4284 133038 4340
rect 133186 4284 133196 4340
rect 133252 4284 137340 4340
rect 137396 4284 137406 4340
rect 141250 4284 141260 4340
rect 141316 4284 143500 4340
rect 143556 4284 143566 4340
rect 147074 4284 147084 4340
rect 147140 4284 148316 4340
rect 148372 4284 148382 4340
rect 163986 4284 163996 4340
rect 164052 4284 165452 4340
rect 165508 4284 165518 4340
rect 49970 4172 49980 4228
rect 50036 4172 50540 4228
rect 50596 4172 57036 4228
rect 57092 4172 57102 4228
rect 120082 4172 120092 4228
rect 120148 4172 137788 4228
rect 140242 4172 140252 4228
rect 140308 4172 143052 4228
rect 143108 4172 144508 4228
rect 144564 4172 144574 4228
rect 147410 4172 147420 4228
rect 147476 4172 153692 4228
rect 153748 4172 154140 4228
rect 154196 4172 154206 4228
rect 165666 4172 165676 4228
rect 165732 4172 184492 4228
rect 184548 4172 184558 4228
rect 57362 4060 57372 4116
rect 57428 4060 58604 4116
rect 58660 4060 58670 4116
rect 68114 4060 68124 4116
rect 68180 4060 69356 4116
rect 69412 4060 69422 4116
rect 103618 4060 103628 4116
rect 103684 4060 130844 4116
rect 130900 4060 130910 4116
rect 132962 4060 132972 4116
rect 133028 4060 133756 4116
rect 133812 4060 133822 4116
rect 137732 4004 137788 4172
rect 137732 3948 149436 4004
rect 149492 3948 150332 4004
rect 150388 3948 150398 4004
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 65906 3892 65916 3948
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 66180 3892 66190 3948
rect 96626 3892 96636 3948
rect 96692 3892 96740 3948
rect 96796 3892 96844 3948
rect 96900 3892 96910 3948
rect 127346 3892 127356 3948
rect 127412 3892 127460 3948
rect 127516 3892 127564 3948
rect 127620 3892 127630 3948
rect 158066 3892 158076 3948
rect 158132 3892 158180 3948
rect 158236 3892 158284 3948
rect 158340 3892 158350 3948
rect 188786 3892 188796 3948
rect 188852 3892 188900 3948
rect 188956 3892 189004 3948
rect 189060 3892 189070 3948
rect 151442 3836 151452 3892
rect 151508 3836 152460 3892
rect 152516 3836 153580 3892
rect 153636 3836 154476 3892
rect 154532 3836 154542 3892
rect 161634 3836 161644 3892
rect 161700 3836 163324 3892
rect 163380 3836 163390 3892
rect 164322 3836 164332 3892
rect 164388 3836 175868 3892
rect 175924 3836 175934 3892
rect 55412 3724 78988 3780
rect 90178 3724 90188 3780
rect 90244 3724 116844 3780
rect 116900 3724 116910 3780
rect 117058 3724 117068 3780
rect 117124 3724 152012 3780
rect 152068 3724 156044 3780
rect 156100 3724 156110 3780
rect 156212 3724 157388 3780
rect 157444 3724 157454 3780
rect 160626 3724 160636 3780
rect 160692 3724 173180 3780
rect 173236 3724 173246 3780
rect 184772 3724 186620 3780
rect 186676 3724 186686 3780
rect 55412 3668 55468 3724
rect 78932 3668 78988 3724
rect 156212 3668 156268 3724
rect 184772 3668 184828 3724
rect 27794 3612 27804 3668
rect 27860 3612 28588 3668
rect 28644 3612 28654 3668
rect 42354 3612 42364 3668
rect 42420 3612 42924 3668
rect 42980 3612 55468 3668
rect 56018 3612 56028 3668
rect 56084 3612 56094 3668
rect 62738 3612 62748 3668
rect 62804 3612 63980 3668
rect 64036 3612 64046 3668
rect 67442 3612 67452 3668
rect 67508 3612 67518 3668
rect 73490 3612 73500 3668
rect 73556 3612 74284 3668
rect 74340 3612 74350 3668
rect 76514 3612 76524 3668
rect 76580 3612 77196 3668
rect 77252 3612 77262 3668
rect 78932 3612 93996 3668
rect 94052 3612 94062 3668
rect 95554 3612 95564 3668
rect 95620 3612 135324 3668
rect 135380 3612 135390 3668
rect 140914 3612 140924 3668
rect 140980 3612 142828 3668
rect 142884 3612 143612 3668
rect 143668 3612 143678 3668
rect 146066 3612 146076 3668
rect 146132 3612 148652 3668
rect 148708 3612 149548 3668
rect 152786 3612 152796 3668
rect 152852 3612 156268 3668
rect 166898 3612 166908 3668
rect 166964 3612 184828 3668
rect 196532 3612 211596 3668
rect 211652 3612 211662 3668
rect 50418 3500 50428 3556
rect 50484 3500 51884 3556
rect 51940 3500 51950 3556
rect 53106 3500 53116 3556
rect 53172 3500 55020 3556
rect 55076 3500 55086 3556
rect 56028 3444 56084 3612
rect 58482 3500 58492 3556
rect 58548 3500 59500 3556
rect 59556 3500 59566 3556
rect 61170 3500 61180 3556
rect 61236 3500 62972 3556
rect 63028 3500 63038 3556
rect 63858 3500 63868 3556
rect 63924 3500 66444 3556
rect 66500 3500 66510 3556
rect 67452 3444 67508 3612
rect 69234 3500 69244 3556
rect 69300 3500 70924 3556
rect 70980 3500 70990 3556
rect 101042 3500 101052 3556
rect 101108 3500 131292 3556
rect 131348 3500 131358 3556
rect 38546 3388 38556 3444
rect 38612 3388 40572 3444
rect 40628 3388 40638 3444
rect 46610 3388 46620 3444
rect 46676 3388 47628 3444
rect 47684 3388 47694 3444
rect 51986 3388 51996 3444
rect 52052 3388 52892 3444
rect 52948 3388 52958 3444
rect 54674 3388 54684 3444
rect 54740 3388 56084 3444
rect 65426 3388 65436 3444
rect 65492 3388 67508 3444
rect 70802 3388 70812 3444
rect 70868 3388 71932 3444
rect 71988 3388 71998 3444
rect 84354 3388 84364 3444
rect 84420 3388 84924 3444
rect 84980 3388 87388 3444
rect 87444 3388 87454 3444
rect 149492 3332 149548 3612
rect 196532 3556 196588 3612
rect 151442 3500 151452 3556
rect 151508 3500 153356 3556
rect 153412 3500 155708 3556
rect 155764 3500 155774 3556
rect 155922 3500 155932 3556
rect 155988 3500 196588 3556
rect 151330 3388 151340 3444
rect 151396 3388 152572 3444
rect 152628 3388 152638 3444
rect 154130 3388 154140 3444
rect 154196 3388 155036 3444
rect 155092 3388 156604 3444
rect 156660 3388 156670 3444
rect 157378 3388 157388 3444
rect 157444 3388 158172 3444
rect 158228 3388 158238 3444
rect 159506 3388 159516 3444
rect 159572 3388 160076 3444
rect 160132 3388 160142 3444
rect 161970 3388 161980 3444
rect 162036 3388 163660 3444
rect 163716 3388 163726 3444
rect 167570 3388 167580 3444
rect 167636 3388 168140 3444
rect 168196 3388 168206 3444
rect 172946 3388 172956 3444
rect 173012 3388 173516 3444
rect 173572 3388 173582 3444
rect 181010 3388 181020 3444
rect 181076 3388 181580 3444
rect 181636 3388 181646 3444
rect 186386 3388 186396 3444
rect 186452 3388 186844 3444
rect 186900 3388 186910 3444
rect 194450 3388 194460 3444
rect 194516 3388 195020 3444
rect 195076 3388 195086 3444
rect 149492 3276 205996 3332
rect 206052 3276 206062 3332
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 50546 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50830 3164
rect 81266 3108 81276 3164
rect 81332 3108 81380 3164
rect 81436 3108 81484 3164
rect 81540 3108 81550 3164
rect 111986 3108 111996 3164
rect 112052 3108 112100 3164
rect 112156 3108 112204 3164
rect 112260 3108 112270 3164
rect 142706 3108 142716 3164
rect 142772 3108 142820 3164
rect 142876 3108 142924 3164
rect 142980 3108 142990 3164
rect 173426 3108 173436 3164
rect 173492 3108 173540 3164
rect 173596 3108 173644 3164
rect 173700 3108 173710 3164
rect 204146 3108 204156 3164
rect 204212 3108 204260 3164
rect 204316 3108 204364 3164
rect 204420 3108 204430 3164
rect 135090 2940 135100 2996
rect 135156 2940 163212 2996
rect 163268 2940 163278 2996
rect 139346 2828 139356 2884
rect 139412 2828 164444 2884
rect 164500 2828 164510 2884
rect 136546 2716 136556 2772
rect 136612 2716 160748 2772
rect 160804 2716 160814 2772
rect 141026 2604 141036 2660
rect 141092 2604 156380 2660
rect 156436 2604 156446 2660
rect 87378 2492 87388 2548
rect 87444 2492 152908 2548
rect 152964 2492 152974 2548
rect 122434 2380 122444 2436
rect 122500 2380 147308 2436
rect 147364 2380 147374 2436
rect 148306 2380 148316 2436
rect 148372 2380 182252 2436
rect 182308 2380 182318 2436
rect 80546 2268 80556 2324
rect 80612 2268 151228 2324
rect 151284 2268 151294 2324
rect 144498 2156 144508 2212
rect 144564 2156 197932 2212
rect 197988 2156 197998 2212
rect 144386 1596 144396 1652
rect 144452 1596 203980 1652
rect 204036 1596 204046 1652
rect 149202 1484 149212 1540
rect 149268 1484 208684 1540
rect 208740 1484 208750 1540
rect 145394 1372 145404 1428
rect 145460 1372 200620 1428
rect 200676 1372 200686 1428
<< via3 >>
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 65916 46228 65972 46284
rect 66020 46228 66076 46284
rect 66124 46228 66180 46284
rect 96636 46228 96692 46284
rect 96740 46228 96796 46284
rect 96844 46228 96900 46284
rect 127356 46228 127412 46284
rect 127460 46228 127516 46284
rect 127564 46228 127620 46284
rect 158076 46228 158132 46284
rect 158180 46228 158236 46284
rect 158284 46228 158340 46284
rect 188796 46228 188852 46284
rect 188900 46228 188956 46284
rect 189004 46228 189060 46284
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 50556 45444 50612 45500
rect 50660 45444 50716 45500
rect 50764 45444 50820 45500
rect 81276 45444 81332 45500
rect 81380 45444 81436 45500
rect 81484 45444 81540 45500
rect 111996 45444 112052 45500
rect 112100 45444 112156 45500
rect 112204 45444 112260 45500
rect 142716 45444 142772 45500
rect 142820 45444 142876 45500
rect 142924 45444 142980 45500
rect 173436 45444 173492 45500
rect 173540 45444 173596 45500
rect 173644 45444 173700 45500
rect 204156 45444 204212 45500
rect 204260 45444 204316 45500
rect 204364 45444 204420 45500
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 65916 44660 65972 44716
rect 66020 44660 66076 44716
rect 66124 44660 66180 44716
rect 96636 44660 96692 44716
rect 96740 44660 96796 44716
rect 96844 44660 96900 44716
rect 127356 44660 127412 44716
rect 127460 44660 127516 44716
rect 127564 44660 127620 44716
rect 158076 44660 158132 44716
rect 158180 44660 158236 44716
rect 158284 44660 158340 44716
rect 188796 44660 188852 44716
rect 188900 44660 188956 44716
rect 189004 44660 189060 44716
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 50556 43876 50612 43932
rect 50660 43876 50716 43932
rect 50764 43876 50820 43932
rect 81276 43876 81332 43932
rect 81380 43876 81436 43932
rect 81484 43876 81540 43932
rect 111996 43876 112052 43932
rect 112100 43876 112156 43932
rect 112204 43876 112260 43932
rect 142716 43876 142772 43932
rect 142820 43876 142876 43932
rect 142924 43876 142980 43932
rect 173436 43876 173492 43932
rect 173540 43876 173596 43932
rect 173644 43876 173700 43932
rect 204156 43876 204212 43932
rect 204260 43876 204316 43932
rect 204364 43876 204420 43932
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 65916 43092 65972 43148
rect 66020 43092 66076 43148
rect 66124 43092 66180 43148
rect 96636 43092 96692 43148
rect 96740 43092 96796 43148
rect 96844 43092 96900 43148
rect 127356 43092 127412 43148
rect 127460 43092 127516 43148
rect 127564 43092 127620 43148
rect 158076 43092 158132 43148
rect 158180 43092 158236 43148
rect 158284 43092 158340 43148
rect 188796 43092 188852 43148
rect 188900 43092 188956 43148
rect 189004 43092 189060 43148
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 50556 42308 50612 42364
rect 50660 42308 50716 42364
rect 50764 42308 50820 42364
rect 81276 42308 81332 42364
rect 81380 42308 81436 42364
rect 81484 42308 81540 42364
rect 111996 42308 112052 42364
rect 112100 42308 112156 42364
rect 112204 42308 112260 42364
rect 142716 42308 142772 42364
rect 142820 42308 142876 42364
rect 142924 42308 142980 42364
rect 173436 42308 173492 42364
rect 173540 42308 173596 42364
rect 173644 42308 173700 42364
rect 204156 42308 204212 42364
rect 204260 42308 204316 42364
rect 204364 42308 204420 42364
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 65916 41524 65972 41580
rect 66020 41524 66076 41580
rect 66124 41524 66180 41580
rect 96636 41524 96692 41580
rect 96740 41524 96796 41580
rect 96844 41524 96900 41580
rect 127356 41524 127412 41580
rect 127460 41524 127516 41580
rect 127564 41524 127620 41580
rect 158076 41524 158132 41580
rect 158180 41524 158236 41580
rect 158284 41524 158340 41580
rect 188796 41524 188852 41580
rect 188900 41524 188956 41580
rect 189004 41524 189060 41580
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 50556 40740 50612 40796
rect 50660 40740 50716 40796
rect 50764 40740 50820 40796
rect 81276 40740 81332 40796
rect 81380 40740 81436 40796
rect 81484 40740 81540 40796
rect 111996 40740 112052 40796
rect 112100 40740 112156 40796
rect 112204 40740 112260 40796
rect 142716 40740 142772 40796
rect 142820 40740 142876 40796
rect 142924 40740 142980 40796
rect 173436 40740 173492 40796
rect 173540 40740 173596 40796
rect 173644 40740 173700 40796
rect 204156 40740 204212 40796
rect 204260 40740 204316 40796
rect 204364 40740 204420 40796
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 65916 39956 65972 40012
rect 66020 39956 66076 40012
rect 66124 39956 66180 40012
rect 96636 39956 96692 40012
rect 96740 39956 96796 40012
rect 96844 39956 96900 40012
rect 127356 39956 127412 40012
rect 127460 39956 127516 40012
rect 127564 39956 127620 40012
rect 158076 39956 158132 40012
rect 158180 39956 158236 40012
rect 158284 39956 158340 40012
rect 188796 39956 188852 40012
rect 188900 39956 188956 40012
rect 189004 39956 189060 40012
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 50556 39172 50612 39228
rect 50660 39172 50716 39228
rect 50764 39172 50820 39228
rect 81276 39172 81332 39228
rect 81380 39172 81436 39228
rect 81484 39172 81540 39228
rect 111996 39172 112052 39228
rect 112100 39172 112156 39228
rect 112204 39172 112260 39228
rect 142716 39172 142772 39228
rect 142820 39172 142876 39228
rect 142924 39172 142980 39228
rect 173436 39172 173492 39228
rect 173540 39172 173596 39228
rect 173644 39172 173700 39228
rect 204156 39172 204212 39228
rect 204260 39172 204316 39228
rect 204364 39172 204420 39228
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 65916 38388 65972 38444
rect 66020 38388 66076 38444
rect 66124 38388 66180 38444
rect 96636 38388 96692 38444
rect 96740 38388 96796 38444
rect 96844 38388 96900 38444
rect 127356 38388 127412 38444
rect 127460 38388 127516 38444
rect 127564 38388 127620 38444
rect 158076 38388 158132 38444
rect 158180 38388 158236 38444
rect 158284 38388 158340 38444
rect 188796 38388 188852 38444
rect 188900 38388 188956 38444
rect 189004 38388 189060 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 50556 37604 50612 37660
rect 50660 37604 50716 37660
rect 50764 37604 50820 37660
rect 81276 37604 81332 37660
rect 81380 37604 81436 37660
rect 81484 37604 81540 37660
rect 111996 37604 112052 37660
rect 112100 37604 112156 37660
rect 112204 37604 112260 37660
rect 142716 37604 142772 37660
rect 142820 37604 142876 37660
rect 142924 37604 142980 37660
rect 173436 37604 173492 37660
rect 173540 37604 173596 37660
rect 173644 37604 173700 37660
rect 204156 37604 204212 37660
rect 204260 37604 204316 37660
rect 204364 37604 204420 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 65916 36820 65972 36876
rect 66020 36820 66076 36876
rect 66124 36820 66180 36876
rect 96636 36820 96692 36876
rect 96740 36820 96796 36876
rect 96844 36820 96900 36876
rect 127356 36820 127412 36876
rect 127460 36820 127516 36876
rect 127564 36820 127620 36876
rect 158076 36820 158132 36876
rect 158180 36820 158236 36876
rect 158284 36820 158340 36876
rect 188796 36820 188852 36876
rect 188900 36820 188956 36876
rect 189004 36820 189060 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 50556 36036 50612 36092
rect 50660 36036 50716 36092
rect 50764 36036 50820 36092
rect 81276 36036 81332 36092
rect 81380 36036 81436 36092
rect 81484 36036 81540 36092
rect 111996 36036 112052 36092
rect 112100 36036 112156 36092
rect 112204 36036 112260 36092
rect 142716 36036 142772 36092
rect 142820 36036 142876 36092
rect 142924 36036 142980 36092
rect 173436 36036 173492 36092
rect 173540 36036 173596 36092
rect 173644 36036 173700 36092
rect 204156 36036 204212 36092
rect 204260 36036 204316 36092
rect 204364 36036 204420 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 65916 35252 65972 35308
rect 66020 35252 66076 35308
rect 66124 35252 66180 35308
rect 96636 35252 96692 35308
rect 96740 35252 96796 35308
rect 96844 35252 96900 35308
rect 127356 35252 127412 35308
rect 127460 35252 127516 35308
rect 127564 35252 127620 35308
rect 158076 35252 158132 35308
rect 158180 35252 158236 35308
rect 158284 35252 158340 35308
rect 188796 35252 188852 35308
rect 188900 35252 188956 35308
rect 189004 35252 189060 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 50556 34468 50612 34524
rect 50660 34468 50716 34524
rect 50764 34468 50820 34524
rect 81276 34468 81332 34524
rect 81380 34468 81436 34524
rect 81484 34468 81540 34524
rect 111996 34468 112052 34524
rect 112100 34468 112156 34524
rect 112204 34468 112260 34524
rect 142716 34468 142772 34524
rect 142820 34468 142876 34524
rect 142924 34468 142980 34524
rect 173436 34468 173492 34524
rect 173540 34468 173596 34524
rect 173644 34468 173700 34524
rect 204156 34468 204212 34524
rect 204260 34468 204316 34524
rect 204364 34468 204420 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 65916 33684 65972 33740
rect 66020 33684 66076 33740
rect 66124 33684 66180 33740
rect 96636 33684 96692 33740
rect 96740 33684 96796 33740
rect 96844 33684 96900 33740
rect 127356 33684 127412 33740
rect 127460 33684 127516 33740
rect 127564 33684 127620 33740
rect 158076 33684 158132 33740
rect 158180 33684 158236 33740
rect 158284 33684 158340 33740
rect 188796 33684 188852 33740
rect 188900 33684 188956 33740
rect 189004 33684 189060 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 50556 32900 50612 32956
rect 50660 32900 50716 32956
rect 50764 32900 50820 32956
rect 81276 32900 81332 32956
rect 81380 32900 81436 32956
rect 81484 32900 81540 32956
rect 111996 32900 112052 32956
rect 112100 32900 112156 32956
rect 112204 32900 112260 32956
rect 142716 32900 142772 32956
rect 142820 32900 142876 32956
rect 142924 32900 142980 32956
rect 173436 32900 173492 32956
rect 173540 32900 173596 32956
rect 173644 32900 173700 32956
rect 204156 32900 204212 32956
rect 204260 32900 204316 32956
rect 204364 32900 204420 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 65916 32116 65972 32172
rect 66020 32116 66076 32172
rect 66124 32116 66180 32172
rect 96636 32116 96692 32172
rect 96740 32116 96796 32172
rect 96844 32116 96900 32172
rect 127356 32116 127412 32172
rect 127460 32116 127516 32172
rect 127564 32116 127620 32172
rect 158076 32116 158132 32172
rect 158180 32116 158236 32172
rect 158284 32116 158340 32172
rect 188796 32116 188852 32172
rect 188900 32116 188956 32172
rect 189004 32116 189060 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 50556 31332 50612 31388
rect 50660 31332 50716 31388
rect 50764 31332 50820 31388
rect 81276 31332 81332 31388
rect 81380 31332 81436 31388
rect 81484 31332 81540 31388
rect 111996 31332 112052 31388
rect 112100 31332 112156 31388
rect 112204 31332 112260 31388
rect 142716 31332 142772 31388
rect 142820 31332 142876 31388
rect 142924 31332 142980 31388
rect 173436 31332 173492 31388
rect 173540 31332 173596 31388
rect 173644 31332 173700 31388
rect 204156 31332 204212 31388
rect 204260 31332 204316 31388
rect 204364 31332 204420 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 65916 30548 65972 30604
rect 66020 30548 66076 30604
rect 66124 30548 66180 30604
rect 96636 30548 96692 30604
rect 96740 30548 96796 30604
rect 96844 30548 96900 30604
rect 127356 30548 127412 30604
rect 127460 30548 127516 30604
rect 127564 30548 127620 30604
rect 158076 30548 158132 30604
rect 158180 30548 158236 30604
rect 158284 30548 158340 30604
rect 188796 30548 188852 30604
rect 188900 30548 188956 30604
rect 189004 30548 189060 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 50556 29764 50612 29820
rect 50660 29764 50716 29820
rect 50764 29764 50820 29820
rect 81276 29764 81332 29820
rect 81380 29764 81436 29820
rect 81484 29764 81540 29820
rect 111996 29764 112052 29820
rect 112100 29764 112156 29820
rect 112204 29764 112260 29820
rect 142716 29764 142772 29820
rect 142820 29764 142876 29820
rect 142924 29764 142980 29820
rect 173436 29764 173492 29820
rect 173540 29764 173596 29820
rect 173644 29764 173700 29820
rect 204156 29764 204212 29820
rect 204260 29764 204316 29820
rect 204364 29764 204420 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 65916 28980 65972 29036
rect 66020 28980 66076 29036
rect 66124 28980 66180 29036
rect 96636 28980 96692 29036
rect 96740 28980 96796 29036
rect 96844 28980 96900 29036
rect 127356 28980 127412 29036
rect 127460 28980 127516 29036
rect 127564 28980 127620 29036
rect 158076 28980 158132 29036
rect 158180 28980 158236 29036
rect 158284 28980 158340 29036
rect 188796 28980 188852 29036
rect 188900 28980 188956 29036
rect 189004 28980 189060 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 50556 28196 50612 28252
rect 50660 28196 50716 28252
rect 50764 28196 50820 28252
rect 81276 28196 81332 28252
rect 81380 28196 81436 28252
rect 81484 28196 81540 28252
rect 111996 28196 112052 28252
rect 112100 28196 112156 28252
rect 112204 28196 112260 28252
rect 142716 28196 142772 28252
rect 142820 28196 142876 28252
rect 142924 28196 142980 28252
rect 173436 28196 173492 28252
rect 173540 28196 173596 28252
rect 173644 28196 173700 28252
rect 204156 28196 204212 28252
rect 204260 28196 204316 28252
rect 204364 28196 204420 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 65916 27412 65972 27468
rect 66020 27412 66076 27468
rect 66124 27412 66180 27468
rect 96636 27412 96692 27468
rect 96740 27412 96796 27468
rect 96844 27412 96900 27468
rect 127356 27412 127412 27468
rect 127460 27412 127516 27468
rect 127564 27412 127620 27468
rect 158076 27412 158132 27468
rect 158180 27412 158236 27468
rect 158284 27412 158340 27468
rect 188796 27412 188852 27468
rect 188900 27412 188956 27468
rect 189004 27412 189060 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 50556 26628 50612 26684
rect 50660 26628 50716 26684
rect 50764 26628 50820 26684
rect 81276 26628 81332 26684
rect 81380 26628 81436 26684
rect 81484 26628 81540 26684
rect 111996 26628 112052 26684
rect 112100 26628 112156 26684
rect 112204 26628 112260 26684
rect 142716 26628 142772 26684
rect 142820 26628 142876 26684
rect 142924 26628 142980 26684
rect 173436 26628 173492 26684
rect 173540 26628 173596 26684
rect 173644 26628 173700 26684
rect 204156 26628 204212 26684
rect 204260 26628 204316 26684
rect 204364 26628 204420 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 65916 25844 65972 25900
rect 66020 25844 66076 25900
rect 66124 25844 66180 25900
rect 96636 25844 96692 25900
rect 96740 25844 96796 25900
rect 96844 25844 96900 25900
rect 127356 25844 127412 25900
rect 127460 25844 127516 25900
rect 127564 25844 127620 25900
rect 158076 25844 158132 25900
rect 158180 25844 158236 25900
rect 158284 25844 158340 25900
rect 188796 25844 188852 25900
rect 188900 25844 188956 25900
rect 189004 25844 189060 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 50556 25060 50612 25116
rect 50660 25060 50716 25116
rect 50764 25060 50820 25116
rect 81276 25060 81332 25116
rect 81380 25060 81436 25116
rect 81484 25060 81540 25116
rect 111996 25060 112052 25116
rect 112100 25060 112156 25116
rect 112204 25060 112260 25116
rect 142716 25060 142772 25116
rect 142820 25060 142876 25116
rect 142924 25060 142980 25116
rect 173436 25060 173492 25116
rect 173540 25060 173596 25116
rect 173644 25060 173700 25116
rect 204156 25060 204212 25116
rect 204260 25060 204316 25116
rect 204364 25060 204420 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 65916 24276 65972 24332
rect 66020 24276 66076 24332
rect 66124 24276 66180 24332
rect 96636 24276 96692 24332
rect 96740 24276 96796 24332
rect 96844 24276 96900 24332
rect 127356 24276 127412 24332
rect 127460 24276 127516 24332
rect 127564 24276 127620 24332
rect 158076 24276 158132 24332
rect 158180 24276 158236 24332
rect 158284 24276 158340 24332
rect 188796 24276 188852 24332
rect 188900 24276 188956 24332
rect 189004 24276 189060 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 50556 23492 50612 23548
rect 50660 23492 50716 23548
rect 50764 23492 50820 23548
rect 81276 23492 81332 23548
rect 81380 23492 81436 23548
rect 81484 23492 81540 23548
rect 111996 23492 112052 23548
rect 112100 23492 112156 23548
rect 112204 23492 112260 23548
rect 142716 23492 142772 23548
rect 142820 23492 142876 23548
rect 142924 23492 142980 23548
rect 173436 23492 173492 23548
rect 173540 23492 173596 23548
rect 173644 23492 173700 23548
rect 204156 23492 204212 23548
rect 204260 23492 204316 23548
rect 204364 23492 204420 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 65916 22708 65972 22764
rect 66020 22708 66076 22764
rect 66124 22708 66180 22764
rect 96636 22708 96692 22764
rect 96740 22708 96796 22764
rect 96844 22708 96900 22764
rect 127356 22708 127412 22764
rect 127460 22708 127516 22764
rect 127564 22708 127620 22764
rect 158076 22708 158132 22764
rect 158180 22708 158236 22764
rect 158284 22708 158340 22764
rect 188796 22708 188852 22764
rect 188900 22708 188956 22764
rect 189004 22708 189060 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 50556 21924 50612 21980
rect 50660 21924 50716 21980
rect 50764 21924 50820 21980
rect 81276 21924 81332 21980
rect 81380 21924 81436 21980
rect 81484 21924 81540 21980
rect 111996 21924 112052 21980
rect 112100 21924 112156 21980
rect 112204 21924 112260 21980
rect 142716 21924 142772 21980
rect 142820 21924 142876 21980
rect 142924 21924 142980 21980
rect 173436 21924 173492 21980
rect 173540 21924 173596 21980
rect 173644 21924 173700 21980
rect 204156 21924 204212 21980
rect 204260 21924 204316 21980
rect 204364 21924 204420 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 65916 21140 65972 21196
rect 66020 21140 66076 21196
rect 66124 21140 66180 21196
rect 96636 21140 96692 21196
rect 96740 21140 96796 21196
rect 96844 21140 96900 21196
rect 127356 21140 127412 21196
rect 127460 21140 127516 21196
rect 127564 21140 127620 21196
rect 158076 21140 158132 21196
rect 158180 21140 158236 21196
rect 158284 21140 158340 21196
rect 188796 21140 188852 21196
rect 188900 21140 188956 21196
rect 189004 21140 189060 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 50556 20356 50612 20412
rect 50660 20356 50716 20412
rect 50764 20356 50820 20412
rect 81276 20356 81332 20412
rect 81380 20356 81436 20412
rect 81484 20356 81540 20412
rect 111996 20356 112052 20412
rect 112100 20356 112156 20412
rect 112204 20356 112260 20412
rect 142716 20356 142772 20412
rect 142820 20356 142876 20412
rect 142924 20356 142980 20412
rect 173436 20356 173492 20412
rect 173540 20356 173596 20412
rect 173644 20356 173700 20412
rect 204156 20356 204212 20412
rect 204260 20356 204316 20412
rect 204364 20356 204420 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 65916 19572 65972 19628
rect 66020 19572 66076 19628
rect 66124 19572 66180 19628
rect 96636 19572 96692 19628
rect 96740 19572 96796 19628
rect 96844 19572 96900 19628
rect 127356 19572 127412 19628
rect 127460 19572 127516 19628
rect 127564 19572 127620 19628
rect 158076 19572 158132 19628
rect 158180 19572 158236 19628
rect 158284 19572 158340 19628
rect 188796 19572 188852 19628
rect 188900 19572 188956 19628
rect 189004 19572 189060 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 50556 18788 50612 18844
rect 50660 18788 50716 18844
rect 50764 18788 50820 18844
rect 81276 18788 81332 18844
rect 81380 18788 81436 18844
rect 81484 18788 81540 18844
rect 111996 18788 112052 18844
rect 112100 18788 112156 18844
rect 112204 18788 112260 18844
rect 142716 18788 142772 18844
rect 142820 18788 142876 18844
rect 142924 18788 142980 18844
rect 173436 18788 173492 18844
rect 173540 18788 173596 18844
rect 173644 18788 173700 18844
rect 204156 18788 204212 18844
rect 204260 18788 204316 18844
rect 204364 18788 204420 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 65916 18004 65972 18060
rect 66020 18004 66076 18060
rect 66124 18004 66180 18060
rect 96636 18004 96692 18060
rect 96740 18004 96796 18060
rect 96844 18004 96900 18060
rect 127356 18004 127412 18060
rect 127460 18004 127516 18060
rect 127564 18004 127620 18060
rect 158076 18004 158132 18060
rect 158180 18004 158236 18060
rect 158284 18004 158340 18060
rect 188796 18004 188852 18060
rect 188900 18004 188956 18060
rect 189004 18004 189060 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 50556 17220 50612 17276
rect 50660 17220 50716 17276
rect 50764 17220 50820 17276
rect 81276 17220 81332 17276
rect 81380 17220 81436 17276
rect 81484 17220 81540 17276
rect 111996 17220 112052 17276
rect 112100 17220 112156 17276
rect 112204 17220 112260 17276
rect 142716 17220 142772 17276
rect 142820 17220 142876 17276
rect 142924 17220 142980 17276
rect 173436 17220 173492 17276
rect 173540 17220 173596 17276
rect 173644 17220 173700 17276
rect 204156 17220 204212 17276
rect 204260 17220 204316 17276
rect 204364 17220 204420 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 65916 16436 65972 16492
rect 66020 16436 66076 16492
rect 66124 16436 66180 16492
rect 96636 16436 96692 16492
rect 96740 16436 96796 16492
rect 96844 16436 96900 16492
rect 127356 16436 127412 16492
rect 127460 16436 127516 16492
rect 127564 16436 127620 16492
rect 158076 16436 158132 16492
rect 158180 16436 158236 16492
rect 158284 16436 158340 16492
rect 188796 16436 188852 16492
rect 188900 16436 188956 16492
rect 189004 16436 189060 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 50556 15652 50612 15708
rect 50660 15652 50716 15708
rect 50764 15652 50820 15708
rect 81276 15652 81332 15708
rect 81380 15652 81436 15708
rect 81484 15652 81540 15708
rect 111996 15652 112052 15708
rect 112100 15652 112156 15708
rect 112204 15652 112260 15708
rect 142716 15652 142772 15708
rect 142820 15652 142876 15708
rect 142924 15652 142980 15708
rect 173436 15652 173492 15708
rect 173540 15652 173596 15708
rect 173644 15652 173700 15708
rect 204156 15652 204212 15708
rect 204260 15652 204316 15708
rect 204364 15652 204420 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 65916 14868 65972 14924
rect 66020 14868 66076 14924
rect 66124 14868 66180 14924
rect 96636 14868 96692 14924
rect 96740 14868 96796 14924
rect 96844 14868 96900 14924
rect 127356 14868 127412 14924
rect 127460 14868 127516 14924
rect 127564 14868 127620 14924
rect 158076 14868 158132 14924
rect 158180 14868 158236 14924
rect 158284 14868 158340 14924
rect 188796 14868 188852 14924
rect 188900 14868 188956 14924
rect 189004 14868 189060 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 50556 14084 50612 14140
rect 50660 14084 50716 14140
rect 50764 14084 50820 14140
rect 81276 14084 81332 14140
rect 81380 14084 81436 14140
rect 81484 14084 81540 14140
rect 111996 14084 112052 14140
rect 112100 14084 112156 14140
rect 112204 14084 112260 14140
rect 142716 14084 142772 14140
rect 142820 14084 142876 14140
rect 142924 14084 142980 14140
rect 173436 14084 173492 14140
rect 173540 14084 173596 14140
rect 173644 14084 173700 14140
rect 204156 14084 204212 14140
rect 204260 14084 204316 14140
rect 204364 14084 204420 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 65916 13300 65972 13356
rect 66020 13300 66076 13356
rect 66124 13300 66180 13356
rect 96636 13300 96692 13356
rect 96740 13300 96796 13356
rect 96844 13300 96900 13356
rect 127356 13300 127412 13356
rect 127460 13300 127516 13356
rect 127564 13300 127620 13356
rect 158076 13300 158132 13356
rect 158180 13300 158236 13356
rect 158284 13300 158340 13356
rect 188796 13300 188852 13356
rect 188900 13300 188956 13356
rect 189004 13300 189060 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 50556 12516 50612 12572
rect 50660 12516 50716 12572
rect 50764 12516 50820 12572
rect 81276 12516 81332 12572
rect 81380 12516 81436 12572
rect 81484 12516 81540 12572
rect 111996 12516 112052 12572
rect 112100 12516 112156 12572
rect 112204 12516 112260 12572
rect 142716 12516 142772 12572
rect 142820 12516 142876 12572
rect 142924 12516 142980 12572
rect 173436 12516 173492 12572
rect 173540 12516 173596 12572
rect 173644 12516 173700 12572
rect 204156 12516 204212 12572
rect 204260 12516 204316 12572
rect 204364 12516 204420 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 65916 11732 65972 11788
rect 66020 11732 66076 11788
rect 66124 11732 66180 11788
rect 96636 11732 96692 11788
rect 96740 11732 96796 11788
rect 96844 11732 96900 11788
rect 127356 11732 127412 11788
rect 127460 11732 127516 11788
rect 127564 11732 127620 11788
rect 158076 11732 158132 11788
rect 158180 11732 158236 11788
rect 158284 11732 158340 11788
rect 188796 11732 188852 11788
rect 188900 11732 188956 11788
rect 189004 11732 189060 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 50556 10948 50612 11004
rect 50660 10948 50716 11004
rect 50764 10948 50820 11004
rect 81276 10948 81332 11004
rect 81380 10948 81436 11004
rect 81484 10948 81540 11004
rect 111996 10948 112052 11004
rect 112100 10948 112156 11004
rect 112204 10948 112260 11004
rect 142716 10948 142772 11004
rect 142820 10948 142876 11004
rect 142924 10948 142980 11004
rect 173436 10948 173492 11004
rect 173540 10948 173596 11004
rect 173644 10948 173700 11004
rect 204156 10948 204212 11004
rect 204260 10948 204316 11004
rect 204364 10948 204420 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 65916 10164 65972 10220
rect 66020 10164 66076 10220
rect 66124 10164 66180 10220
rect 96636 10164 96692 10220
rect 96740 10164 96796 10220
rect 96844 10164 96900 10220
rect 127356 10164 127412 10220
rect 127460 10164 127516 10220
rect 127564 10164 127620 10220
rect 158076 10164 158132 10220
rect 158180 10164 158236 10220
rect 158284 10164 158340 10220
rect 188796 10164 188852 10220
rect 188900 10164 188956 10220
rect 189004 10164 189060 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 50556 9380 50612 9436
rect 50660 9380 50716 9436
rect 50764 9380 50820 9436
rect 81276 9380 81332 9436
rect 81380 9380 81436 9436
rect 81484 9380 81540 9436
rect 111996 9380 112052 9436
rect 112100 9380 112156 9436
rect 112204 9380 112260 9436
rect 142716 9380 142772 9436
rect 142820 9380 142876 9436
rect 142924 9380 142980 9436
rect 173436 9380 173492 9436
rect 173540 9380 173596 9436
rect 173644 9380 173700 9436
rect 204156 9380 204212 9436
rect 204260 9380 204316 9436
rect 204364 9380 204420 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 65916 8596 65972 8652
rect 66020 8596 66076 8652
rect 66124 8596 66180 8652
rect 96636 8596 96692 8652
rect 96740 8596 96796 8652
rect 96844 8596 96900 8652
rect 127356 8596 127412 8652
rect 127460 8596 127516 8652
rect 127564 8596 127620 8652
rect 158076 8596 158132 8652
rect 158180 8596 158236 8652
rect 158284 8596 158340 8652
rect 188796 8596 188852 8652
rect 188900 8596 188956 8652
rect 189004 8596 189060 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 50556 7812 50612 7868
rect 50660 7812 50716 7868
rect 50764 7812 50820 7868
rect 81276 7812 81332 7868
rect 81380 7812 81436 7868
rect 81484 7812 81540 7868
rect 111996 7812 112052 7868
rect 112100 7812 112156 7868
rect 112204 7812 112260 7868
rect 142716 7812 142772 7868
rect 142820 7812 142876 7868
rect 142924 7812 142980 7868
rect 173436 7812 173492 7868
rect 173540 7812 173596 7868
rect 173644 7812 173700 7868
rect 204156 7812 204212 7868
rect 204260 7812 204316 7868
rect 204364 7812 204420 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 65916 7028 65972 7084
rect 66020 7028 66076 7084
rect 66124 7028 66180 7084
rect 96636 7028 96692 7084
rect 96740 7028 96796 7084
rect 96844 7028 96900 7084
rect 127356 7028 127412 7084
rect 127460 7028 127516 7084
rect 127564 7028 127620 7084
rect 158076 7028 158132 7084
rect 158180 7028 158236 7084
rect 158284 7028 158340 7084
rect 188796 7028 188852 7084
rect 188900 7028 188956 7084
rect 189004 7028 189060 7084
rect 162764 6972 162820 7028
rect 163996 6412 164052 6468
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 50556 6244 50612 6300
rect 50660 6244 50716 6300
rect 50764 6244 50820 6300
rect 81276 6244 81332 6300
rect 81380 6244 81436 6300
rect 81484 6244 81540 6300
rect 111996 6244 112052 6300
rect 112100 6244 112156 6300
rect 112204 6244 112260 6300
rect 142716 6244 142772 6300
rect 142820 6244 142876 6300
rect 142924 6244 142980 6300
rect 173436 6244 173492 6300
rect 173540 6244 173596 6300
rect 173644 6244 173700 6300
rect 204156 6244 204212 6300
rect 204260 6244 204316 6300
rect 204364 6244 204420 6300
rect 162764 6076 162820 6132
rect 163548 6076 163604 6132
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 65916 5460 65972 5516
rect 66020 5460 66076 5516
rect 66124 5460 66180 5516
rect 96636 5460 96692 5516
rect 96740 5460 96796 5516
rect 96844 5460 96900 5516
rect 127356 5460 127412 5516
rect 127460 5460 127516 5516
rect 127564 5460 127620 5516
rect 158076 5460 158132 5516
rect 158180 5460 158236 5516
rect 158284 5460 158340 5516
rect 188796 5460 188852 5516
rect 188900 5460 188956 5516
rect 189004 5460 189060 5516
rect 163996 5180 164052 5236
rect 163548 4844 163604 4900
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 50556 4676 50612 4732
rect 50660 4676 50716 4732
rect 50764 4676 50820 4732
rect 81276 4676 81332 4732
rect 81380 4676 81436 4732
rect 81484 4676 81540 4732
rect 111996 4676 112052 4732
rect 112100 4676 112156 4732
rect 112204 4676 112260 4732
rect 142716 4676 142772 4732
rect 142820 4676 142876 4732
rect 142924 4676 142980 4732
rect 137788 4620 137844 4676
rect 173436 4676 173492 4732
rect 173540 4676 173596 4732
rect 173644 4676 173700 4732
rect 204156 4676 204212 4732
rect 204260 4676 204316 4732
rect 204364 4676 204420 4732
rect 137788 4396 137844 4452
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 65916 3892 65972 3948
rect 66020 3892 66076 3948
rect 66124 3892 66180 3948
rect 96636 3892 96692 3948
rect 96740 3892 96796 3948
rect 96844 3892 96900 3948
rect 127356 3892 127412 3948
rect 127460 3892 127516 3948
rect 127564 3892 127620 3948
rect 158076 3892 158132 3948
rect 158180 3892 158236 3948
rect 158284 3892 158340 3948
rect 188796 3892 188852 3948
rect 188900 3892 188956 3948
rect 189004 3892 189060 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
rect 50556 3108 50612 3164
rect 50660 3108 50716 3164
rect 50764 3108 50820 3164
rect 81276 3108 81332 3164
rect 81380 3108 81436 3164
rect 81484 3108 81540 3164
rect 111996 3108 112052 3164
rect 112100 3108 112156 3164
rect 112204 3108 112260 3164
rect 142716 3108 142772 3164
rect 142820 3108 142876 3164
rect 142924 3108 142980 3164
rect 173436 3108 173492 3164
rect 173540 3108 173596 3164
rect 173644 3108 173700 3164
rect 204156 3108 204212 3164
rect 204260 3108 204316 3164
rect 204364 3108 204420 3164
<< metal4 >>
rect 4448 46284 4768 46316
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 4448 44716 4768 46228
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 45500 20128 46316
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 46284 35488 46316
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
rect 50528 45500 50848 46316
rect 50528 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50848 45500
rect 50528 43932 50848 45444
rect 50528 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50848 43932
rect 50528 42364 50848 43876
rect 50528 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50848 42364
rect 50528 40796 50848 42308
rect 50528 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50848 40796
rect 50528 39228 50848 40740
rect 50528 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50848 39228
rect 50528 37660 50848 39172
rect 50528 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50848 37660
rect 50528 36092 50848 37604
rect 50528 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50848 36092
rect 50528 34524 50848 36036
rect 50528 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50848 34524
rect 50528 32956 50848 34468
rect 50528 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50848 32956
rect 50528 31388 50848 32900
rect 50528 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50848 31388
rect 50528 29820 50848 31332
rect 50528 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50848 29820
rect 50528 28252 50848 29764
rect 50528 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50848 28252
rect 50528 26684 50848 28196
rect 50528 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50848 26684
rect 50528 25116 50848 26628
rect 50528 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50848 25116
rect 50528 23548 50848 25060
rect 50528 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50848 23548
rect 50528 21980 50848 23492
rect 50528 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50848 21980
rect 50528 20412 50848 21924
rect 50528 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50848 20412
rect 50528 18844 50848 20356
rect 50528 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50848 18844
rect 50528 17276 50848 18788
rect 50528 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50848 17276
rect 50528 15708 50848 17220
rect 50528 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50848 15708
rect 50528 14140 50848 15652
rect 50528 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50848 14140
rect 50528 12572 50848 14084
rect 50528 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50848 12572
rect 50528 11004 50848 12516
rect 50528 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50848 11004
rect 50528 9436 50848 10948
rect 50528 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50848 9436
rect 50528 7868 50848 9380
rect 50528 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50848 7868
rect 50528 6300 50848 7812
rect 50528 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50848 6300
rect 50528 4732 50848 6244
rect 50528 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50848 4732
rect 50528 3164 50848 4676
rect 50528 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50848 3164
rect 50528 3076 50848 3108
rect 65888 46284 66208 46316
rect 65888 46228 65916 46284
rect 65972 46228 66020 46284
rect 66076 46228 66124 46284
rect 66180 46228 66208 46284
rect 65888 44716 66208 46228
rect 65888 44660 65916 44716
rect 65972 44660 66020 44716
rect 66076 44660 66124 44716
rect 66180 44660 66208 44716
rect 65888 43148 66208 44660
rect 65888 43092 65916 43148
rect 65972 43092 66020 43148
rect 66076 43092 66124 43148
rect 66180 43092 66208 43148
rect 65888 41580 66208 43092
rect 65888 41524 65916 41580
rect 65972 41524 66020 41580
rect 66076 41524 66124 41580
rect 66180 41524 66208 41580
rect 65888 40012 66208 41524
rect 65888 39956 65916 40012
rect 65972 39956 66020 40012
rect 66076 39956 66124 40012
rect 66180 39956 66208 40012
rect 65888 38444 66208 39956
rect 65888 38388 65916 38444
rect 65972 38388 66020 38444
rect 66076 38388 66124 38444
rect 66180 38388 66208 38444
rect 65888 36876 66208 38388
rect 65888 36820 65916 36876
rect 65972 36820 66020 36876
rect 66076 36820 66124 36876
rect 66180 36820 66208 36876
rect 65888 35308 66208 36820
rect 65888 35252 65916 35308
rect 65972 35252 66020 35308
rect 66076 35252 66124 35308
rect 66180 35252 66208 35308
rect 65888 33740 66208 35252
rect 65888 33684 65916 33740
rect 65972 33684 66020 33740
rect 66076 33684 66124 33740
rect 66180 33684 66208 33740
rect 65888 32172 66208 33684
rect 65888 32116 65916 32172
rect 65972 32116 66020 32172
rect 66076 32116 66124 32172
rect 66180 32116 66208 32172
rect 65888 30604 66208 32116
rect 65888 30548 65916 30604
rect 65972 30548 66020 30604
rect 66076 30548 66124 30604
rect 66180 30548 66208 30604
rect 65888 29036 66208 30548
rect 65888 28980 65916 29036
rect 65972 28980 66020 29036
rect 66076 28980 66124 29036
rect 66180 28980 66208 29036
rect 65888 27468 66208 28980
rect 65888 27412 65916 27468
rect 65972 27412 66020 27468
rect 66076 27412 66124 27468
rect 66180 27412 66208 27468
rect 65888 25900 66208 27412
rect 65888 25844 65916 25900
rect 65972 25844 66020 25900
rect 66076 25844 66124 25900
rect 66180 25844 66208 25900
rect 65888 24332 66208 25844
rect 65888 24276 65916 24332
rect 65972 24276 66020 24332
rect 66076 24276 66124 24332
rect 66180 24276 66208 24332
rect 65888 22764 66208 24276
rect 65888 22708 65916 22764
rect 65972 22708 66020 22764
rect 66076 22708 66124 22764
rect 66180 22708 66208 22764
rect 65888 21196 66208 22708
rect 65888 21140 65916 21196
rect 65972 21140 66020 21196
rect 66076 21140 66124 21196
rect 66180 21140 66208 21196
rect 65888 19628 66208 21140
rect 65888 19572 65916 19628
rect 65972 19572 66020 19628
rect 66076 19572 66124 19628
rect 66180 19572 66208 19628
rect 65888 18060 66208 19572
rect 65888 18004 65916 18060
rect 65972 18004 66020 18060
rect 66076 18004 66124 18060
rect 66180 18004 66208 18060
rect 65888 16492 66208 18004
rect 65888 16436 65916 16492
rect 65972 16436 66020 16492
rect 66076 16436 66124 16492
rect 66180 16436 66208 16492
rect 65888 14924 66208 16436
rect 65888 14868 65916 14924
rect 65972 14868 66020 14924
rect 66076 14868 66124 14924
rect 66180 14868 66208 14924
rect 65888 13356 66208 14868
rect 65888 13300 65916 13356
rect 65972 13300 66020 13356
rect 66076 13300 66124 13356
rect 66180 13300 66208 13356
rect 65888 11788 66208 13300
rect 65888 11732 65916 11788
rect 65972 11732 66020 11788
rect 66076 11732 66124 11788
rect 66180 11732 66208 11788
rect 65888 10220 66208 11732
rect 65888 10164 65916 10220
rect 65972 10164 66020 10220
rect 66076 10164 66124 10220
rect 66180 10164 66208 10220
rect 65888 8652 66208 10164
rect 65888 8596 65916 8652
rect 65972 8596 66020 8652
rect 66076 8596 66124 8652
rect 66180 8596 66208 8652
rect 65888 7084 66208 8596
rect 65888 7028 65916 7084
rect 65972 7028 66020 7084
rect 66076 7028 66124 7084
rect 66180 7028 66208 7084
rect 65888 5516 66208 7028
rect 65888 5460 65916 5516
rect 65972 5460 66020 5516
rect 66076 5460 66124 5516
rect 66180 5460 66208 5516
rect 65888 3948 66208 5460
rect 65888 3892 65916 3948
rect 65972 3892 66020 3948
rect 66076 3892 66124 3948
rect 66180 3892 66208 3948
rect 65888 3076 66208 3892
rect 81248 45500 81568 46316
rect 81248 45444 81276 45500
rect 81332 45444 81380 45500
rect 81436 45444 81484 45500
rect 81540 45444 81568 45500
rect 81248 43932 81568 45444
rect 81248 43876 81276 43932
rect 81332 43876 81380 43932
rect 81436 43876 81484 43932
rect 81540 43876 81568 43932
rect 81248 42364 81568 43876
rect 81248 42308 81276 42364
rect 81332 42308 81380 42364
rect 81436 42308 81484 42364
rect 81540 42308 81568 42364
rect 81248 40796 81568 42308
rect 81248 40740 81276 40796
rect 81332 40740 81380 40796
rect 81436 40740 81484 40796
rect 81540 40740 81568 40796
rect 81248 39228 81568 40740
rect 81248 39172 81276 39228
rect 81332 39172 81380 39228
rect 81436 39172 81484 39228
rect 81540 39172 81568 39228
rect 81248 37660 81568 39172
rect 81248 37604 81276 37660
rect 81332 37604 81380 37660
rect 81436 37604 81484 37660
rect 81540 37604 81568 37660
rect 81248 36092 81568 37604
rect 81248 36036 81276 36092
rect 81332 36036 81380 36092
rect 81436 36036 81484 36092
rect 81540 36036 81568 36092
rect 81248 34524 81568 36036
rect 81248 34468 81276 34524
rect 81332 34468 81380 34524
rect 81436 34468 81484 34524
rect 81540 34468 81568 34524
rect 81248 32956 81568 34468
rect 81248 32900 81276 32956
rect 81332 32900 81380 32956
rect 81436 32900 81484 32956
rect 81540 32900 81568 32956
rect 81248 31388 81568 32900
rect 81248 31332 81276 31388
rect 81332 31332 81380 31388
rect 81436 31332 81484 31388
rect 81540 31332 81568 31388
rect 81248 29820 81568 31332
rect 81248 29764 81276 29820
rect 81332 29764 81380 29820
rect 81436 29764 81484 29820
rect 81540 29764 81568 29820
rect 81248 28252 81568 29764
rect 81248 28196 81276 28252
rect 81332 28196 81380 28252
rect 81436 28196 81484 28252
rect 81540 28196 81568 28252
rect 81248 26684 81568 28196
rect 81248 26628 81276 26684
rect 81332 26628 81380 26684
rect 81436 26628 81484 26684
rect 81540 26628 81568 26684
rect 81248 25116 81568 26628
rect 81248 25060 81276 25116
rect 81332 25060 81380 25116
rect 81436 25060 81484 25116
rect 81540 25060 81568 25116
rect 81248 23548 81568 25060
rect 81248 23492 81276 23548
rect 81332 23492 81380 23548
rect 81436 23492 81484 23548
rect 81540 23492 81568 23548
rect 81248 21980 81568 23492
rect 81248 21924 81276 21980
rect 81332 21924 81380 21980
rect 81436 21924 81484 21980
rect 81540 21924 81568 21980
rect 81248 20412 81568 21924
rect 81248 20356 81276 20412
rect 81332 20356 81380 20412
rect 81436 20356 81484 20412
rect 81540 20356 81568 20412
rect 81248 18844 81568 20356
rect 81248 18788 81276 18844
rect 81332 18788 81380 18844
rect 81436 18788 81484 18844
rect 81540 18788 81568 18844
rect 81248 17276 81568 18788
rect 81248 17220 81276 17276
rect 81332 17220 81380 17276
rect 81436 17220 81484 17276
rect 81540 17220 81568 17276
rect 81248 15708 81568 17220
rect 81248 15652 81276 15708
rect 81332 15652 81380 15708
rect 81436 15652 81484 15708
rect 81540 15652 81568 15708
rect 81248 14140 81568 15652
rect 81248 14084 81276 14140
rect 81332 14084 81380 14140
rect 81436 14084 81484 14140
rect 81540 14084 81568 14140
rect 81248 12572 81568 14084
rect 81248 12516 81276 12572
rect 81332 12516 81380 12572
rect 81436 12516 81484 12572
rect 81540 12516 81568 12572
rect 81248 11004 81568 12516
rect 81248 10948 81276 11004
rect 81332 10948 81380 11004
rect 81436 10948 81484 11004
rect 81540 10948 81568 11004
rect 81248 9436 81568 10948
rect 81248 9380 81276 9436
rect 81332 9380 81380 9436
rect 81436 9380 81484 9436
rect 81540 9380 81568 9436
rect 81248 7868 81568 9380
rect 81248 7812 81276 7868
rect 81332 7812 81380 7868
rect 81436 7812 81484 7868
rect 81540 7812 81568 7868
rect 81248 6300 81568 7812
rect 81248 6244 81276 6300
rect 81332 6244 81380 6300
rect 81436 6244 81484 6300
rect 81540 6244 81568 6300
rect 81248 4732 81568 6244
rect 81248 4676 81276 4732
rect 81332 4676 81380 4732
rect 81436 4676 81484 4732
rect 81540 4676 81568 4732
rect 81248 3164 81568 4676
rect 81248 3108 81276 3164
rect 81332 3108 81380 3164
rect 81436 3108 81484 3164
rect 81540 3108 81568 3164
rect 81248 3076 81568 3108
rect 96608 46284 96928 46316
rect 96608 46228 96636 46284
rect 96692 46228 96740 46284
rect 96796 46228 96844 46284
rect 96900 46228 96928 46284
rect 96608 44716 96928 46228
rect 96608 44660 96636 44716
rect 96692 44660 96740 44716
rect 96796 44660 96844 44716
rect 96900 44660 96928 44716
rect 96608 43148 96928 44660
rect 96608 43092 96636 43148
rect 96692 43092 96740 43148
rect 96796 43092 96844 43148
rect 96900 43092 96928 43148
rect 96608 41580 96928 43092
rect 96608 41524 96636 41580
rect 96692 41524 96740 41580
rect 96796 41524 96844 41580
rect 96900 41524 96928 41580
rect 96608 40012 96928 41524
rect 96608 39956 96636 40012
rect 96692 39956 96740 40012
rect 96796 39956 96844 40012
rect 96900 39956 96928 40012
rect 96608 38444 96928 39956
rect 96608 38388 96636 38444
rect 96692 38388 96740 38444
rect 96796 38388 96844 38444
rect 96900 38388 96928 38444
rect 96608 36876 96928 38388
rect 96608 36820 96636 36876
rect 96692 36820 96740 36876
rect 96796 36820 96844 36876
rect 96900 36820 96928 36876
rect 96608 35308 96928 36820
rect 96608 35252 96636 35308
rect 96692 35252 96740 35308
rect 96796 35252 96844 35308
rect 96900 35252 96928 35308
rect 96608 33740 96928 35252
rect 96608 33684 96636 33740
rect 96692 33684 96740 33740
rect 96796 33684 96844 33740
rect 96900 33684 96928 33740
rect 96608 32172 96928 33684
rect 96608 32116 96636 32172
rect 96692 32116 96740 32172
rect 96796 32116 96844 32172
rect 96900 32116 96928 32172
rect 96608 30604 96928 32116
rect 96608 30548 96636 30604
rect 96692 30548 96740 30604
rect 96796 30548 96844 30604
rect 96900 30548 96928 30604
rect 96608 29036 96928 30548
rect 96608 28980 96636 29036
rect 96692 28980 96740 29036
rect 96796 28980 96844 29036
rect 96900 28980 96928 29036
rect 96608 27468 96928 28980
rect 96608 27412 96636 27468
rect 96692 27412 96740 27468
rect 96796 27412 96844 27468
rect 96900 27412 96928 27468
rect 96608 25900 96928 27412
rect 96608 25844 96636 25900
rect 96692 25844 96740 25900
rect 96796 25844 96844 25900
rect 96900 25844 96928 25900
rect 96608 24332 96928 25844
rect 96608 24276 96636 24332
rect 96692 24276 96740 24332
rect 96796 24276 96844 24332
rect 96900 24276 96928 24332
rect 96608 22764 96928 24276
rect 96608 22708 96636 22764
rect 96692 22708 96740 22764
rect 96796 22708 96844 22764
rect 96900 22708 96928 22764
rect 96608 21196 96928 22708
rect 96608 21140 96636 21196
rect 96692 21140 96740 21196
rect 96796 21140 96844 21196
rect 96900 21140 96928 21196
rect 96608 19628 96928 21140
rect 96608 19572 96636 19628
rect 96692 19572 96740 19628
rect 96796 19572 96844 19628
rect 96900 19572 96928 19628
rect 96608 18060 96928 19572
rect 96608 18004 96636 18060
rect 96692 18004 96740 18060
rect 96796 18004 96844 18060
rect 96900 18004 96928 18060
rect 96608 16492 96928 18004
rect 96608 16436 96636 16492
rect 96692 16436 96740 16492
rect 96796 16436 96844 16492
rect 96900 16436 96928 16492
rect 96608 14924 96928 16436
rect 96608 14868 96636 14924
rect 96692 14868 96740 14924
rect 96796 14868 96844 14924
rect 96900 14868 96928 14924
rect 96608 13356 96928 14868
rect 96608 13300 96636 13356
rect 96692 13300 96740 13356
rect 96796 13300 96844 13356
rect 96900 13300 96928 13356
rect 96608 11788 96928 13300
rect 96608 11732 96636 11788
rect 96692 11732 96740 11788
rect 96796 11732 96844 11788
rect 96900 11732 96928 11788
rect 96608 10220 96928 11732
rect 96608 10164 96636 10220
rect 96692 10164 96740 10220
rect 96796 10164 96844 10220
rect 96900 10164 96928 10220
rect 96608 8652 96928 10164
rect 96608 8596 96636 8652
rect 96692 8596 96740 8652
rect 96796 8596 96844 8652
rect 96900 8596 96928 8652
rect 96608 7084 96928 8596
rect 96608 7028 96636 7084
rect 96692 7028 96740 7084
rect 96796 7028 96844 7084
rect 96900 7028 96928 7084
rect 96608 5516 96928 7028
rect 96608 5460 96636 5516
rect 96692 5460 96740 5516
rect 96796 5460 96844 5516
rect 96900 5460 96928 5516
rect 96608 3948 96928 5460
rect 96608 3892 96636 3948
rect 96692 3892 96740 3948
rect 96796 3892 96844 3948
rect 96900 3892 96928 3948
rect 96608 3076 96928 3892
rect 111968 45500 112288 46316
rect 111968 45444 111996 45500
rect 112052 45444 112100 45500
rect 112156 45444 112204 45500
rect 112260 45444 112288 45500
rect 111968 43932 112288 45444
rect 111968 43876 111996 43932
rect 112052 43876 112100 43932
rect 112156 43876 112204 43932
rect 112260 43876 112288 43932
rect 111968 42364 112288 43876
rect 111968 42308 111996 42364
rect 112052 42308 112100 42364
rect 112156 42308 112204 42364
rect 112260 42308 112288 42364
rect 111968 40796 112288 42308
rect 111968 40740 111996 40796
rect 112052 40740 112100 40796
rect 112156 40740 112204 40796
rect 112260 40740 112288 40796
rect 111968 39228 112288 40740
rect 111968 39172 111996 39228
rect 112052 39172 112100 39228
rect 112156 39172 112204 39228
rect 112260 39172 112288 39228
rect 111968 37660 112288 39172
rect 111968 37604 111996 37660
rect 112052 37604 112100 37660
rect 112156 37604 112204 37660
rect 112260 37604 112288 37660
rect 111968 36092 112288 37604
rect 111968 36036 111996 36092
rect 112052 36036 112100 36092
rect 112156 36036 112204 36092
rect 112260 36036 112288 36092
rect 111968 34524 112288 36036
rect 111968 34468 111996 34524
rect 112052 34468 112100 34524
rect 112156 34468 112204 34524
rect 112260 34468 112288 34524
rect 111968 32956 112288 34468
rect 111968 32900 111996 32956
rect 112052 32900 112100 32956
rect 112156 32900 112204 32956
rect 112260 32900 112288 32956
rect 111968 31388 112288 32900
rect 111968 31332 111996 31388
rect 112052 31332 112100 31388
rect 112156 31332 112204 31388
rect 112260 31332 112288 31388
rect 111968 29820 112288 31332
rect 111968 29764 111996 29820
rect 112052 29764 112100 29820
rect 112156 29764 112204 29820
rect 112260 29764 112288 29820
rect 111968 28252 112288 29764
rect 111968 28196 111996 28252
rect 112052 28196 112100 28252
rect 112156 28196 112204 28252
rect 112260 28196 112288 28252
rect 111968 26684 112288 28196
rect 111968 26628 111996 26684
rect 112052 26628 112100 26684
rect 112156 26628 112204 26684
rect 112260 26628 112288 26684
rect 111968 25116 112288 26628
rect 111968 25060 111996 25116
rect 112052 25060 112100 25116
rect 112156 25060 112204 25116
rect 112260 25060 112288 25116
rect 111968 23548 112288 25060
rect 111968 23492 111996 23548
rect 112052 23492 112100 23548
rect 112156 23492 112204 23548
rect 112260 23492 112288 23548
rect 111968 21980 112288 23492
rect 111968 21924 111996 21980
rect 112052 21924 112100 21980
rect 112156 21924 112204 21980
rect 112260 21924 112288 21980
rect 111968 20412 112288 21924
rect 111968 20356 111996 20412
rect 112052 20356 112100 20412
rect 112156 20356 112204 20412
rect 112260 20356 112288 20412
rect 111968 18844 112288 20356
rect 111968 18788 111996 18844
rect 112052 18788 112100 18844
rect 112156 18788 112204 18844
rect 112260 18788 112288 18844
rect 111968 17276 112288 18788
rect 111968 17220 111996 17276
rect 112052 17220 112100 17276
rect 112156 17220 112204 17276
rect 112260 17220 112288 17276
rect 111968 15708 112288 17220
rect 111968 15652 111996 15708
rect 112052 15652 112100 15708
rect 112156 15652 112204 15708
rect 112260 15652 112288 15708
rect 111968 14140 112288 15652
rect 111968 14084 111996 14140
rect 112052 14084 112100 14140
rect 112156 14084 112204 14140
rect 112260 14084 112288 14140
rect 111968 12572 112288 14084
rect 111968 12516 111996 12572
rect 112052 12516 112100 12572
rect 112156 12516 112204 12572
rect 112260 12516 112288 12572
rect 111968 11004 112288 12516
rect 111968 10948 111996 11004
rect 112052 10948 112100 11004
rect 112156 10948 112204 11004
rect 112260 10948 112288 11004
rect 111968 9436 112288 10948
rect 111968 9380 111996 9436
rect 112052 9380 112100 9436
rect 112156 9380 112204 9436
rect 112260 9380 112288 9436
rect 111968 7868 112288 9380
rect 111968 7812 111996 7868
rect 112052 7812 112100 7868
rect 112156 7812 112204 7868
rect 112260 7812 112288 7868
rect 111968 6300 112288 7812
rect 111968 6244 111996 6300
rect 112052 6244 112100 6300
rect 112156 6244 112204 6300
rect 112260 6244 112288 6300
rect 111968 4732 112288 6244
rect 111968 4676 111996 4732
rect 112052 4676 112100 4732
rect 112156 4676 112204 4732
rect 112260 4676 112288 4732
rect 111968 3164 112288 4676
rect 111968 3108 111996 3164
rect 112052 3108 112100 3164
rect 112156 3108 112204 3164
rect 112260 3108 112288 3164
rect 111968 3076 112288 3108
rect 127328 46284 127648 46316
rect 127328 46228 127356 46284
rect 127412 46228 127460 46284
rect 127516 46228 127564 46284
rect 127620 46228 127648 46284
rect 127328 44716 127648 46228
rect 127328 44660 127356 44716
rect 127412 44660 127460 44716
rect 127516 44660 127564 44716
rect 127620 44660 127648 44716
rect 127328 43148 127648 44660
rect 127328 43092 127356 43148
rect 127412 43092 127460 43148
rect 127516 43092 127564 43148
rect 127620 43092 127648 43148
rect 127328 41580 127648 43092
rect 127328 41524 127356 41580
rect 127412 41524 127460 41580
rect 127516 41524 127564 41580
rect 127620 41524 127648 41580
rect 127328 40012 127648 41524
rect 127328 39956 127356 40012
rect 127412 39956 127460 40012
rect 127516 39956 127564 40012
rect 127620 39956 127648 40012
rect 127328 38444 127648 39956
rect 127328 38388 127356 38444
rect 127412 38388 127460 38444
rect 127516 38388 127564 38444
rect 127620 38388 127648 38444
rect 127328 36876 127648 38388
rect 127328 36820 127356 36876
rect 127412 36820 127460 36876
rect 127516 36820 127564 36876
rect 127620 36820 127648 36876
rect 127328 35308 127648 36820
rect 127328 35252 127356 35308
rect 127412 35252 127460 35308
rect 127516 35252 127564 35308
rect 127620 35252 127648 35308
rect 127328 33740 127648 35252
rect 127328 33684 127356 33740
rect 127412 33684 127460 33740
rect 127516 33684 127564 33740
rect 127620 33684 127648 33740
rect 127328 32172 127648 33684
rect 127328 32116 127356 32172
rect 127412 32116 127460 32172
rect 127516 32116 127564 32172
rect 127620 32116 127648 32172
rect 127328 30604 127648 32116
rect 127328 30548 127356 30604
rect 127412 30548 127460 30604
rect 127516 30548 127564 30604
rect 127620 30548 127648 30604
rect 127328 29036 127648 30548
rect 127328 28980 127356 29036
rect 127412 28980 127460 29036
rect 127516 28980 127564 29036
rect 127620 28980 127648 29036
rect 127328 27468 127648 28980
rect 127328 27412 127356 27468
rect 127412 27412 127460 27468
rect 127516 27412 127564 27468
rect 127620 27412 127648 27468
rect 127328 25900 127648 27412
rect 127328 25844 127356 25900
rect 127412 25844 127460 25900
rect 127516 25844 127564 25900
rect 127620 25844 127648 25900
rect 127328 24332 127648 25844
rect 127328 24276 127356 24332
rect 127412 24276 127460 24332
rect 127516 24276 127564 24332
rect 127620 24276 127648 24332
rect 127328 22764 127648 24276
rect 127328 22708 127356 22764
rect 127412 22708 127460 22764
rect 127516 22708 127564 22764
rect 127620 22708 127648 22764
rect 127328 21196 127648 22708
rect 127328 21140 127356 21196
rect 127412 21140 127460 21196
rect 127516 21140 127564 21196
rect 127620 21140 127648 21196
rect 127328 19628 127648 21140
rect 127328 19572 127356 19628
rect 127412 19572 127460 19628
rect 127516 19572 127564 19628
rect 127620 19572 127648 19628
rect 127328 18060 127648 19572
rect 127328 18004 127356 18060
rect 127412 18004 127460 18060
rect 127516 18004 127564 18060
rect 127620 18004 127648 18060
rect 127328 16492 127648 18004
rect 127328 16436 127356 16492
rect 127412 16436 127460 16492
rect 127516 16436 127564 16492
rect 127620 16436 127648 16492
rect 127328 14924 127648 16436
rect 127328 14868 127356 14924
rect 127412 14868 127460 14924
rect 127516 14868 127564 14924
rect 127620 14868 127648 14924
rect 127328 13356 127648 14868
rect 127328 13300 127356 13356
rect 127412 13300 127460 13356
rect 127516 13300 127564 13356
rect 127620 13300 127648 13356
rect 127328 11788 127648 13300
rect 127328 11732 127356 11788
rect 127412 11732 127460 11788
rect 127516 11732 127564 11788
rect 127620 11732 127648 11788
rect 127328 10220 127648 11732
rect 127328 10164 127356 10220
rect 127412 10164 127460 10220
rect 127516 10164 127564 10220
rect 127620 10164 127648 10220
rect 127328 8652 127648 10164
rect 127328 8596 127356 8652
rect 127412 8596 127460 8652
rect 127516 8596 127564 8652
rect 127620 8596 127648 8652
rect 127328 7084 127648 8596
rect 127328 7028 127356 7084
rect 127412 7028 127460 7084
rect 127516 7028 127564 7084
rect 127620 7028 127648 7084
rect 127328 5516 127648 7028
rect 127328 5460 127356 5516
rect 127412 5460 127460 5516
rect 127516 5460 127564 5516
rect 127620 5460 127648 5516
rect 127328 3948 127648 5460
rect 142688 45500 143008 46316
rect 142688 45444 142716 45500
rect 142772 45444 142820 45500
rect 142876 45444 142924 45500
rect 142980 45444 143008 45500
rect 142688 43932 143008 45444
rect 142688 43876 142716 43932
rect 142772 43876 142820 43932
rect 142876 43876 142924 43932
rect 142980 43876 143008 43932
rect 142688 42364 143008 43876
rect 142688 42308 142716 42364
rect 142772 42308 142820 42364
rect 142876 42308 142924 42364
rect 142980 42308 143008 42364
rect 142688 40796 143008 42308
rect 142688 40740 142716 40796
rect 142772 40740 142820 40796
rect 142876 40740 142924 40796
rect 142980 40740 143008 40796
rect 142688 39228 143008 40740
rect 142688 39172 142716 39228
rect 142772 39172 142820 39228
rect 142876 39172 142924 39228
rect 142980 39172 143008 39228
rect 142688 37660 143008 39172
rect 142688 37604 142716 37660
rect 142772 37604 142820 37660
rect 142876 37604 142924 37660
rect 142980 37604 143008 37660
rect 142688 36092 143008 37604
rect 142688 36036 142716 36092
rect 142772 36036 142820 36092
rect 142876 36036 142924 36092
rect 142980 36036 143008 36092
rect 142688 34524 143008 36036
rect 142688 34468 142716 34524
rect 142772 34468 142820 34524
rect 142876 34468 142924 34524
rect 142980 34468 143008 34524
rect 142688 32956 143008 34468
rect 142688 32900 142716 32956
rect 142772 32900 142820 32956
rect 142876 32900 142924 32956
rect 142980 32900 143008 32956
rect 142688 31388 143008 32900
rect 142688 31332 142716 31388
rect 142772 31332 142820 31388
rect 142876 31332 142924 31388
rect 142980 31332 143008 31388
rect 142688 29820 143008 31332
rect 142688 29764 142716 29820
rect 142772 29764 142820 29820
rect 142876 29764 142924 29820
rect 142980 29764 143008 29820
rect 142688 28252 143008 29764
rect 142688 28196 142716 28252
rect 142772 28196 142820 28252
rect 142876 28196 142924 28252
rect 142980 28196 143008 28252
rect 142688 26684 143008 28196
rect 142688 26628 142716 26684
rect 142772 26628 142820 26684
rect 142876 26628 142924 26684
rect 142980 26628 143008 26684
rect 142688 25116 143008 26628
rect 142688 25060 142716 25116
rect 142772 25060 142820 25116
rect 142876 25060 142924 25116
rect 142980 25060 143008 25116
rect 142688 23548 143008 25060
rect 142688 23492 142716 23548
rect 142772 23492 142820 23548
rect 142876 23492 142924 23548
rect 142980 23492 143008 23548
rect 142688 21980 143008 23492
rect 142688 21924 142716 21980
rect 142772 21924 142820 21980
rect 142876 21924 142924 21980
rect 142980 21924 143008 21980
rect 142688 20412 143008 21924
rect 142688 20356 142716 20412
rect 142772 20356 142820 20412
rect 142876 20356 142924 20412
rect 142980 20356 143008 20412
rect 142688 18844 143008 20356
rect 142688 18788 142716 18844
rect 142772 18788 142820 18844
rect 142876 18788 142924 18844
rect 142980 18788 143008 18844
rect 142688 17276 143008 18788
rect 142688 17220 142716 17276
rect 142772 17220 142820 17276
rect 142876 17220 142924 17276
rect 142980 17220 143008 17276
rect 142688 15708 143008 17220
rect 142688 15652 142716 15708
rect 142772 15652 142820 15708
rect 142876 15652 142924 15708
rect 142980 15652 143008 15708
rect 142688 14140 143008 15652
rect 142688 14084 142716 14140
rect 142772 14084 142820 14140
rect 142876 14084 142924 14140
rect 142980 14084 143008 14140
rect 142688 12572 143008 14084
rect 142688 12516 142716 12572
rect 142772 12516 142820 12572
rect 142876 12516 142924 12572
rect 142980 12516 143008 12572
rect 142688 11004 143008 12516
rect 142688 10948 142716 11004
rect 142772 10948 142820 11004
rect 142876 10948 142924 11004
rect 142980 10948 143008 11004
rect 142688 9436 143008 10948
rect 142688 9380 142716 9436
rect 142772 9380 142820 9436
rect 142876 9380 142924 9436
rect 142980 9380 143008 9436
rect 142688 7868 143008 9380
rect 142688 7812 142716 7868
rect 142772 7812 142820 7868
rect 142876 7812 142924 7868
rect 142980 7812 143008 7868
rect 142688 6300 143008 7812
rect 142688 6244 142716 6300
rect 142772 6244 142820 6300
rect 142876 6244 142924 6300
rect 142980 6244 143008 6300
rect 142688 4732 143008 6244
rect 137788 4676 137844 4686
rect 137788 4452 137844 4620
rect 137788 4386 137844 4396
rect 142688 4676 142716 4732
rect 142772 4676 142820 4732
rect 142876 4676 142924 4732
rect 142980 4676 143008 4732
rect 127328 3892 127356 3948
rect 127412 3892 127460 3948
rect 127516 3892 127564 3948
rect 127620 3892 127648 3948
rect 127328 3076 127648 3892
rect 142688 3164 143008 4676
rect 142688 3108 142716 3164
rect 142772 3108 142820 3164
rect 142876 3108 142924 3164
rect 142980 3108 143008 3164
rect 142688 3076 143008 3108
rect 158048 46284 158368 46316
rect 158048 46228 158076 46284
rect 158132 46228 158180 46284
rect 158236 46228 158284 46284
rect 158340 46228 158368 46284
rect 158048 44716 158368 46228
rect 158048 44660 158076 44716
rect 158132 44660 158180 44716
rect 158236 44660 158284 44716
rect 158340 44660 158368 44716
rect 158048 43148 158368 44660
rect 158048 43092 158076 43148
rect 158132 43092 158180 43148
rect 158236 43092 158284 43148
rect 158340 43092 158368 43148
rect 158048 41580 158368 43092
rect 158048 41524 158076 41580
rect 158132 41524 158180 41580
rect 158236 41524 158284 41580
rect 158340 41524 158368 41580
rect 158048 40012 158368 41524
rect 158048 39956 158076 40012
rect 158132 39956 158180 40012
rect 158236 39956 158284 40012
rect 158340 39956 158368 40012
rect 158048 38444 158368 39956
rect 158048 38388 158076 38444
rect 158132 38388 158180 38444
rect 158236 38388 158284 38444
rect 158340 38388 158368 38444
rect 158048 36876 158368 38388
rect 158048 36820 158076 36876
rect 158132 36820 158180 36876
rect 158236 36820 158284 36876
rect 158340 36820 158368 36876
rect 158048 35308 158368 36820
rect 158048 35252 158076 35308
rect 158132 35252 158180 35308
rect 158236 35252 158284 35308
rect 158340 35252 158368 35308
rect 158048 33740 158368 35252
rect 158048 33684 158076 33740
rect 158132 33684 158180 33740
rect 158236 33684 158284 33740
rect 158340 33684 158368 33740
rect 158048 32172 158368 33684
rect 158048 32116 158076 32172
rect 158132 32116 158180 32172
rect 158236 32116 158284 32172
rect 158340 32116 158368 32172
rect 158048 30604 158368 32116
rect 158048 30548 158076 30604
rect 158132 30548 158180 30604
rect 158236 30548 158284 30604
rect 158340 30548 158368 30604
rect 158048 29036 158368 30548
rect 158048 28980 158076 29036
rect 158132 28980 158180 29036
rect 158236 28980 158284 29036
rect 158340 28980 158368 29036
rect 158048 27468 158368 28980
rect 158048 27412 158076 27468
rect 158132 27412 158180 27468
rect 158236 27412 158284 27468
rect 158340 27412 158368 27468
rect 158048 25900 158368 27412
rect 158048 25844 158076 25900
rect 158132 25844 158180 25900
rect 158236 25844 158284 25900
rect 158340 25844 158368 25900
rect 158048 24332 158368 25844
rect 158048 24276 158076 24332
rect 158132 24276 158180 24332
rect 158236 24276 158284 24332
rect 158340 24276 158368 24332
rect 158048 22764 158368 24276
rect 158048 22708 158076 22764
rect 158132 22708 158180 22764
rect 158236 22708 158284 22764
rect 158340 22708 158368 22764
rect 158048 21196 158368 22708
rect 158048 21140 158076 21196
rect 158132 21140 158180 21196
rect 158236 21140 158284 21196
rect 158340 21140 158368 21196
rect 158048 19628 158368 21140
rect 158048 19572 158076 19628
rect 158132 19572 158180 19628
rect 158236 19572 158284 19628
rect 158340 19572 158368 19628
rect 158048 18060 158368 19572
rect 158048 18004 158076 18060
rect 158132 18004 158180 18060
rect 158236 18004 158284 18060
rect 158340 18004 158368 18060
rect 158048 16492 158368 18004
rect 158048 16436 158076 16492
rect 158132 16436 158180 16492
rect 158236 16436 158284 16492
rect 158340 16436 158368 16492
rect 158048 14924 158368 16436
rect 158048 14868 158076 14924
rect 158132 14868 158180 14924
rect 158236 14868 158284 14924
rect 158340 14868 158368 14924
rect 158048 13356 158368 14868
rect 158048 13300 158076 13356
rect 158132 13300 158180 13356
rect 158236 13300 158284 13356
rect 158340 13300 158368 13356
rect 158048 11788 158368 13300
rect 158048 11732 158076 11788
rect 158132 11732 158180 11788
rect 158236 11732 158284 11788
rect 158340 11732 158368 11788
rect 158048 10220 158368 11732
rect 158048 10164 158076 10220
rect 158132 10164 158180 10220
rect 158236 10164 158284 10220
rect 158340 10164 158368 10220
rect 158048 8652 158368 10164
rect 158048 8596 158076 8652
rect 158132 8596 158180 8652
rect 158236 8596 158284 8652
rect 158340 8596 158368 8652
rect 158048 7084 158368 8596
rect 158048 7028 158076 7084
rect 158132 7028 158180 7084
rect 158236 7028 158284 7084
rect 158340 7028 158368 7084
rect 173408 45500 173728 46316
rect 173408 45444 173436 45500
rect 173492 45444 173540 45500
rect 173596 45444 173644 45500
rect 173700 45444 173728 45500
rect 173408 43932 173728 45444
rect 173408 43876 173436 43932
rect 173492 43876 173540 43932
rect 173596 43876 173644 43932
rect 173700 43876 173728 43932
rect 173408 42364 173728 43876
rect 173408 42308 173436 42364
rect 173492 42308 173540 42364
rect 173596 42308 173644 42364
rect 173700 42308 173728 42364
rect 173408 40796 173728 42308
rect 173408 40740 173436 40796
rect 173492 40740 173540 40796
rect 173596 40740 173644 40796
rect 173700 40740 173728 40796
rect 173408 39228 173728 40740
rect 173408 39172 173436 39228
rect 173492 39172 173540 39228
rect 173596 39172 173644 39228
rect 173700 39172 173728 39228
rect 173408 37660 173728 39172
rect 173408 37604 173436 37660
rect 173492 37604 173540 37660
rect 173596 37604 173644 37660
rect 173700 37604 173728 37660
rect 173408 36092 173728 37604
rect 173408 36036 173436 36092
rect 173492 36036 173540 36092
rect 173596 36036 173644 36092
rect 173700 36036 173728 36092
rect 173408 34524 173728 36036
rect 173408 34468 173436 34524
rect 173492 34468 173540 34524
rect 173596 34468 173644 34524
rect 173700 34468 173728 34524
rect 173408 32956 173728 34468
rect 173408 32900 173436 32956
rect 173492 32900 173540 32956
rect 173596 32900 173644 32956
rect 173700 32900 173728 32956
rect 173408 31388 173728 32900
rect 173408 31332 173436 31388
rect 173492 31332 173540 31388
rect 173596 31332 173644 31388
rect 173700 31332 173728 31388
rect 173408 29820 173728 31332
rect 173408 29764 173436 29820
rect 173492 29764 173540 29820
rect 173596 29764 173644 29820
rect 173700 29764 173728 29820
rect 173408 28252 173728 29764
rect 173408 28196 173436 28252
rect 173492 28196 173540 28252
rect 173596 28196 173644 28252
rect 173700 28196 173728 28252
rect 173408 26684 173728 28196
rect 173408 26628 173436 26684
rect 173492 26628 173540 26684
rect 173596 26628 173644 26684
rect 173700 26628 173728 26684
rect 173408 25116 173728 26628
rect 173408 25060 173436 25116
rect 173492 25060 173540 25116
rect 173596 25060 173644 25116
rect 173700 25060 173728 25116
rect 173408 23548 173728 25060
rect 173408 23492 173436 23548
rect 173492 23492 173540 23548
rect 173596 23492 173644 23548
rect 173700 23492 173728 23548
rect 173408 21980 173728 23492
rect 173408 21924 173436 21980
rect 173492 21924 173540 21980
rect 173596 21924 173644 21980
rect 173700 21924 173728 21980
rect 173408 20412 173728 21924
rect 173408 20356 173436 20412
rect 173492 20356 173540 20412
rect 173596 20356 173644 20412
rect 173700 20356 173728 20412
rect 173408 18844 173728 20356
rect 173408 18788 173436 18844
rect 173492 18788 173540 18844
rect 173596 18788 173644 18844
rect 173700 18788 173728 18844
rect 173408 17276 173728 18788
rect 173408 17220 173436 17276
rect 173492 17220 173540 17276
rect 173596 17220 173644 17276
rect 173700 17220 173728 17276
rect 173408 15708 173728 17220
rect 173408 15652 173436 15708
rect 173492 15652 173540 15708
rect 173596 15652 173644 15708
rect 173700 15652 173728 15708
rect 173408 14140 173728 15652
rect 173408 14084 173436 14140
rect 173492 14084 173540 14140
rect 173596 14084 173644 14140
rect 173700 14084 173728 14140
rect 173408 12572 173728 14084
rect 173408 12516 173436 12572
rect 173492 12516 173540 12572
rect 173596 12516 173644 12572
rect 173700 12516 173728 12572
rect 173408 11004 173728 12516
rect 173408 10948 173436 11004
rect 173492 10948 173540 11004
rect 173596 10948 173644 11004
rect 173700 10948 173728 11004
rect 173408 9436 173728 10948
rect 173408 9380 173436 9436
rect 173492 9380 173540 9436
rect 173596 9380 173644 9436
rect 173700 9380 173728 9436
rect 173408 7868 173728 9380
rect 173408 7812 173436 7868
rect 173492 7812 173540 7868
rect 173596 7812 173644 7868
rect 173700 7812 173728 7868
rect 158048 5516 158368 7028
rect 162764 7028 162820 7038
rect 162764 6132 162820 6972
rect 163996 6468 164052 6478
rect 162764 6066 162820 6076
rect 163548 6132 163604 6142
rect 158048 5460 158076 5516
rect 158132 5460 158180 5516
rect 158236 5460 158284 5516
rect 158340 5460 158368 5516
rect 158048 3948 158368 5460
rect 163548 4900 163604 6076
rect 163996 5236 164052 6412
rect 163996 5170 164052 5180
rect 173408 6300 173728 7812
rect 173408 6244 173436 6300
rect 173492 6244 173540 6300
rect 173596 6244 173644 6300
rect 173700 6244 173728 6300
rect 163548 4834 163604 4844
rect 158048 3892 158076 3948
rect 158132 3892 158180 3948
rect 158236 3892 158284 3948
rect 158340 3892 158368 3948
rect 158048 3076 158368 3892
rect 173408 4732 173728 6244
rect 173408 4676 173436 4732
rect 173492 4676 173540 4732
rect 173596 4676 173644 4732
rect 173700 4676 173728 4732
rect 173408 3164 173728 4676
rect 173408 3108 173436 3164
rect 173492 3108 173540 3164
rect 173596 3108 173644 3164
rect 173700 3108 173728 3164
rect 173408 3076 173728 3108
rect 188768 46284 189088 46316
rect 188768 46228 188796 46284
rect 188852 46228 188900 46284
rect 188956 46228 189004 46284
rect 189060 46228 189088 46284
rect 188768 44716 189088 46228
rect 188768 44660 188796 44716
rect 188852 44660 188900 44716
rect 188956 44660 189004 44716
rect 189060 44660 189088 44716
rect 188768 43148 189088 44660
rect 188768 43092 188796 43148
rect 188852 43092 188900 43148
rect 188956 43092 189004 43148
rect 189060 43092 189088 43148
rect 188768 41580 189088 43092
rect 188768 41524 188796 41580
rect 188852 41524 188900 41580
rect 188956 41524 189004 41580
rect 189060 41524 189088 41580
rect 188768 40012 189088 41524
rect 188768 39956 188796 40012
rect 188852 39956 188900 40012
rect 188956 39956 189004 40012
rect 189060 39956 189088 40012
rect 188768 38444 189088 39956
rect 188768 38388 188796 38444
rect 188852 38388 188900 38444
rect 188956 38388 189004 38444
rect 189060 38388 189088 38444
rect 188768 36876 189088 38388
rect 188768 36820 188796 36876
rect 188852 36820 188900 36876
rect 188956 36820 189004 36876
rect 189060 36820 189088 36876
rect 188768 35308 189088 36820
rect 188768 35252 188796 35308
rect 188852 35252 188900 35308
rect 188956 35252 189004 35308
rect 189060 35252 189088 35308
rect 188768 33740 189088 35252
rect 188768 33684 188796 33740
rect 188852 33684 188900 33740
rect 188956 33684 189004 33740
rect 189060 33684 189088 33740
rect 188768 32172 189088 33684
rect 188768 32116 188796 32172
rect 188852 32116 188900 32172
rect 188956 32116 189004 32172
rect 189060 32116 189088 32172
rect 188768 30604 189088 32116
rect 188768 30548 188796 30604
rect 188852 30548 188900 30604
rect 188956 30548 189004 30604
rect 189060 30548 189088 30604
rect 188768 29036 189088 30548
rect 188768 28980 188796 29036
rect 188852 28980 188900 29036
rect 188956 28980 189004 29036
rect 189060 28980 189088 29036
rect 188768 27468 189088 28980
rect 188768 27412 188796 27468
rect 188852 27412 188900 27468
rect 188956 27412 189004 27468
rect 189060 27412 189088 27468
rect 188768 25900 189088 27412
rect 188768 25844 188796 25900
rect 188852 25844 188900 25900
rect 188956 25844 189004 25900
rect 189060 25844 189088 25900
rect 188768 24332 189088 25844
rect 188768 24276 188796 24332
rect 188852 24276 188900 24332
rect 188956 24276 189004 24332
rect 189060 24276 189088 24332
rect 188768 22764 189088 24276
rect 188768 22708 188796 22764
rect 188852 22708 188900 22764
rect 188956 22708 189004 22764
rect 189060 22708 189088 22764
rect 188768 21196 189088 22708
rect 188768 21140 188796 21196
rect 188852 21140 188900 21196
rect 188956 21140 189004 21196
rect 189060 21140 189088 21196
rect 188768 19628 189088 21140
rect 188768 19572 188796 19628
rect 188852 19572 188900 19628
rect 188956 19572 189004 19628
rect 189060 19572 189088 19628
rect 188768 18060 189088 19572
rect 188768 18004 188796 18060
rect 188852 18004 188900 18060
rect 188956 18004 189004 18060
rect 189060 18004 189088 18060
rect 188768 16492 189088 18004
rect 188768 16436 188796 16492
rect 188852 16436 188900 16492
rect 188956 16436 189004 16492
rect 189060 16436 189088 16492
rect 188768 14924 189088 16436
rect 188768 14868 188796 14924
rect 188852 14868 188900 14924
rect 188956 14868 189004 14924
rect 189060 14868 189088 14924
rect 188768 13356 189088 14868
rect 188768 13300 188796 13356
rect 188852 13300 188900 13356
rect 188956 13300 189004 13356
rect 189060 13300 189088 13356
rect 188768 11788 189088 13300
rect 188768 11732 188796 11788
rect 188852 11732 188900 11788
rect 188956 11732 189004 11788
rect 189060 11732 189088 11788
rect 188768 10220 189088 11732
rect 188768 10164 188796 10220
rect 188852 10164 188900 10220
rect 188956 10164 189004 10220
rect 189060 10164 189088 10220
rect 188768 8652 189088 10164
rect 188768 8596 188796 8652
rect 188852 8596 188900 8652
rect 188956 8596 189004 8652
rect 189060 8596 189088 8652
rect 188768 7084 189088 8596
rect 188768 7028 188796 7084
rect 188852 7028 188900 7084
rect 188956 7028 189004 7084
rect 189060 7028 189088 7084
rect 188768 5516 189088 7028
rect 188768 5460 188796 5516
rect 188852 5460 188900 5516
rect 188956 5460 189004 5516
rect 189060 5460 189088 5516
rect 188768 3948 189088 5460
rect 188768 3892 188796 3948
rect 188852 3892 188900 3948
rect 188956 3892 189004 3948
rect 189060 3892 189088 3948
rect 188768 3076 189088 3892
rect 204128 45500 204448 46316
rect 204128 45444 204156 45500
rect 204212 45444 204260 45500
rect 204316 45444 204364 45500
rect 204420 45444 204448 45500
rect 204128 43932 204448 45444
rect 204128 43876 204156 43932
rect 204212 43876 204260 43932
rect 204316 43876 204364 43932
rect 204420 43876 204448 43932
rect 204128 42364 204448 43876
rect 204128 42308 204156 42364
rect 204212 42308 204260 42364
rect 204316 42308 204364 42364
rect 204420 42308 204448 42364
rect 204128 40796 204448 42308
rect 204128 40740 204156 40796
rect 204212 40740 204260 40796
rect 204316 40740 204364 40796
rect 204420 40740 204448 40796
rect 204128 39228 204448 40740
rect 204128 39172 204156 39228
rect 204212 39172 204260 39228
rect 204316 39172 204364 39228
rect 204420 39172 204448 39228
rect 204128 37660 204448 39172
rect 204128 37604 204156 37660
rect 204212 37604 204260 37660
rect 204316 37604 204364 37660
rect 204420 37604 204448 37660
rect 204128 36092 204448 37604
rect 204128 36036 204156 36092
rect 204212 36036 204260 36092
rect 204316 36036 204364 36092
rect 204420 36036 204448 36092
rect 204128 34524 204448 36036
rect 204128 34468 204156 34524
rect 204212 34468 204260 34524
rect 204316 34468 204364 34524
rect 204420 34468 204448 34524
rect 204128 32956 204448 34468
rect 204128 32900 204156 32956
rect 204212 32900 204260 32956
rect 204316 32900 204364 32956
rect 204420 32900 204448 32956
rect 204128 31388 204448 32900
rect 204128 31332 204156 31388
rect 204212 31332 204260 31388
rect 204316 31332 204364 31388
rect 204420 31332 204448 31388
rect 204128 29820 204448 31332
rect 204128 29764 204156 29820
rect 204212 29764 204260 29820
rect 204316 29764 204364 29820
rect 204420 29764 204448 29820
rect 204128 28252 204448 29764
rect 204128 28196 204156 28252
rect 204212 28196 204260 28252
rect 204316 28196 204364 28252
rect 204420 28196 204448 28252
rect 204128 26684 204448 28196
rect 204128 26628 204156 26684
rect 204212 26628 204260 26684
rect 204316 26628 204364 26684
rect 204420 26628 204448 26684
rect 204128 25116 204448 26628
rect 204128 25060 204156 25116
rect 204212 25060 204260 25116
rect 204316 25060 204364 25116
rect 204420 25060 204448 25116
rect 204128 23548 204448 25060
rect 204128 23492 204156 23548
rect 204212 23492 204260 23548
rect 204316 23492 204364 23548
rect 204420 23492 204448 23548
rect 204128 21980 204448 23492
rect 204128 21924 204156 21980
rect 204212 21924 204260 21980
rect 204316 21924 204364 21980
rect 204420 21924 204448 21980
rect 204128 20412 204448 21924
rect 204128 20356 204156 20412
rect 204212 20356 204260 20412
rect 204316 20356 204364 20412
rect 204420 20356 204448 20412
rect 204128 18844 204448 20356
rect 204128 18788 204156 18844
rect 204212 18788 204260 18844
rect 204316 18788 204364 18844
rect 204420 18788 204448 18844
rect 204128 17276 204448 18788
rect 204128 17220 204156 17276
rect 204212 17220 204260 17276
rect 204316 17220 204364 17276
rect 204420 17220 204448 17276
rect 204128 15708 204448 17220
rect 204128 15652 204156 15708
rect 204212 15652 204260 15708
rect 204316 15652 204364 15708
rect 204420 15652 204448 15708
rect 204128 14140 204448 15652
rect 204128 14084 204156 14140
rect 204212 14084 204260 14140
rect 204316 14084 204364 14140
rect 204420 14084 204448 14140
rect 204128 12572 204448 14084
rect 204128 12516 204156 12572
rect 204212 12516 204260 12572
rect 204316 12516 204364 12572
rect 204420 12516 204448 12572
rect 204128 11004 204448 12516
rect 204128 10948 204156 11004
rect 204212 10948 204260 11004
rect 204316 10948 204364 11004
rect 204420 10948 204448 11004
rect 204128 9436 204448 10948
rect 204128 9380 204156 9436
rect 204212 9380 204260 9436
rect 204316 9380 204364 9436
rect 204420 9380 204448 9436
rect 204128 7868 204448 9380
rect 204128 7812 204156 7868
rect 204212 7812 204260 7868
rect 204316 7812 204364 7868
rect 204420 7812 204448 7868
rect 204128 6300 204448 7812
rect 204128 6244 204156 6300
rect 204212 6244 204260 6300
rect 204316 6244 204364 6300
rect 204420 6244 204448 6300
rect 204128 4732 204448 6244
rect 204128 4676 204156 4732
rect 204212 4676 204260 4732
rect 204316 4676 204364 4732
rect 204420 4676 204448 4732
rect 204128 3164 204448 4676
rect 204128 3108 204156 3164
rect 204212 3108 204260 3164
rect 204316 3108 204364 3164
rect 204420 3108 204448 3164
rect 204128 3076 204448 3108
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _106_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 161392 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _107_
timestamp 1698431365
transform 1 0 161056 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _108_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 164304 0 1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _109_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 162176 0 -1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _110_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 134624 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _111_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 131488 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _112_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 148736 0 -1 6272
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _113_
timestamp 1698431365
transform 1 0 149296 0 -1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _114_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 164416 0 -1 4704
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _115_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 166544 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _116_
timestamp 1698431365
transform -1 0 164192 0 -1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _117_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 162064 0 1 4704
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _118_
timestamp 1698431365
transform -1 0 135968 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _119_
timestamp 1698431365
transform 1 0 131040 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _120_
timestamp 1698431365
transform -1 0 151872 0 1 4704
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _121_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 151088 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _122_
timestamp 1698431365
transform 1 0 162960 0 -1 7840
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _123_
timestamp 1698431365
transform -1 0 164752 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _124_
timestamp 1698431365
transform -1 0 163296 0 1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_2  _125_
timestamp 1698431365
transform 1 0 163296 0 1 4704
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _126_
timestamp 1698431365
transform -1 0 135968 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _127_
timestamp 1698431365
transform 1 0 131936 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _128_
timestamp 1698431365
transform 1 0 144480 0 -1 7840
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _129_
timestamp 1698431365
transform -1 0 152880 0 1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _130_
timestamp 1698431365
transform 1 0 162176 0 -1 7840
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _131_
timestamp 1698431365
transform 1 0 162512 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _132_
timestamp 1698431365
transform 1 0 161728 0 -1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _133_
timestamp 1698431365
transform -1 0 163520 0 -1 6272
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _134_
timestamp 1698431365
transform -1 0 138432 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _135_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 109872 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _136_
timestamp 1698431365
transform 1 0 148512 0 1 6272
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _137_
timestamp 1698431365
transform 1 0 150528 0 -1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _138_
timestamp 1698431365
transform 1 0 160160 0 1 6272
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _139_
timestamp 1698431365
transform -1 0 161840 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _140_
timestamp 1698431365
transform -1 0 160944 0 -1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _141_
timestamp 1698431365
transform -1 0 161056 0 -1 6272
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _142_
timestamp 1698431365
transform -1 0 138432 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _143_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 137536 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _144_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 136416 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _145_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 141792 0 -1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _146_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 139776 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _147_
timestamp 1698431365
transform 1 0 148960 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _148_
timestamp 1698431365
transform 1 0 151088 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _149_
timestamp 1698431365
transform 1 0 148064 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _150_
timestamp 1698431365
transform 1 0 151760 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _151_
timestamp 1698431365
transform 1 0 148064 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _152_
timestamp 1698431365
transform 1 0 152992 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _153_
timestamp 1698431365
transform -1 0 154112 0 -1 9408
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _154_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 135968 0 1 6272
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _155_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 137200 0 1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _156_
timestamp 1698431365
transform -1 0 148736 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _157_
timestamp 1698431365
transform 1 0 150640 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _158_
timestamp 1698431365
transform 1 0 153888 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _159_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 148400 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _160_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 147840 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _161_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 156688 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _162_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 140560 0 1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _163_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 154784 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _164_
timestamp 1698431365
transform -1 0 151760 0 1 9408
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _165_
timestamp 1698431365
transform -1 0 145600 0 1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _166_
timestamp 1698431365
transform -1 0 140336 0 -1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _167_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 147168 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _168_
timestamp 1698431365
transform 1 0 156688 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _169_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 155792 0 -1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _170_
timestamp 1698431365
transform -1 0 155904 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _171_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 148736 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _172_
timestamp 1698431365
transform 1 0 161056 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_4  _173_
timestamp 1698431365
transform -1 0 157472 0 1 6272
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _174_
timestamp 1698431365
transform 1 0 149968 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _175_
timestamp 1698431365
transform -1 0 151872 0 1 7840
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _176_
timestamp 1698431365
transform -1 0 142016 0 -1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _177_
timestamp 1698431365
transform -1 0 138320 0 1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _178_
timestamp 1698431365
transform 1 0 155904 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _179_
timestamp 1698431365
transform -1 0 156688 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _180_
timestamp 1698431365
transform 1 0 154224 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _181_
timestamp 1698431365
transform -1 0 148960 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  _182_
timestamp 1698431365
transform -1 0 144256 0 -1 7840
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _183_
timestamp 1698431365
transform 1 0 140112 0 -1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _184_
timestamp 1698431365
transform 1 0 133504 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _185_
timestamp 1698431365
transform -1 0 142464 0 -1 4704
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _186_
timestamp 1698431365
transform 1 0 150528 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _187_
timestamp 1698431365
transform -1 0 160832 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _188_
timestamp 1698431365
transform -1 0 153552 0 -1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _189_
timestamp 1698431365
transform -1 0 156016 0 -1 4704
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _190_
timestamp 1698431365
transform 1 0 159152 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _191_
timestamp 1698431365
transform -1 0 164416 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _192_
timestamp 1698431365
transform -1 0 157696 0 1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _193_
timestamp 1698431365
transform -1 0 154224 0 1 4704
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _194_
timestamp 1698431365
transform -1 0 142016 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _195_
timestamp 1698431365
transform 1 0 133952 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _196_
timestamp 1698431365
transform -1 0 144032 0 1 4704
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _197_
timestamp 1698431365
transform 1 0 151536 0 -1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _198_
timestamp 1698431365
transform 1 0 154448 0 1 4704
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _199_
timestamp 1698431365
transform -1 0 163184 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _200_
timestamp 1698431365
transform 1 0 155344 0 1 9408
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _201_
timestamp 1698431365
transform 1 0 155232 0 1 4704
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _202_
timestamp 1698431365
transform -1 0 142352 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _203_
timestamp 1698431365
transform 1 0 135520 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _204_
timestamp 1698431365
transform -1 0 144032 0 1 6272
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _205_
timestamp 1698431365
transform -1 0 152544 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _206_
timestamp 1698431365
transform 1 0 151872 0 1 3136
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _207_
timestamp 1698431365
transform 1 0 156016 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _208_
timestamp 1698431365
transform 1 0 157696 0 1 4704
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _209_
timestamp 1698431365
transform 1 0 162288 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _210_
timestamp 1698431365
transform -1 0 165312 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _211_
timestamp 1698431365
transform 1 0 154672 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _212_
timestamp 1698431365
transform -1 0 157360 0 1 10976
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _213_
timestamp 1698431365
transform -1 0 157696 0 1 4704
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_4  _214_
timestamp 1698431365
transform -1 0 139328 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _215_
timestamp 1698431365
transform 1 0 130256 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _216_
timestamp 1698431365
transform -1 0 135520 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _217_
timestamp 1698431365
transform -1 0 145376 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _218_
timestamp 1698431365
transform 1 0 144032 0 1 4704
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  _219_
timestamp 1698431365
transform -1 0 144256 0 1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_4  _220_
timestamp 1698431365
transform -1 0 148624 0 -1 4704
box -86 -86 5350 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _221_
timestamp 1698431365
transform -1 0 151200 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _222_
timestamp 1698431365
transform 1 0 148624 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _223_
timestamp 1698431365
transform 1 0 149296 0 -1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _224_
timestamp 1698431365
transform 1 0 161280 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _225_
timestamp 1698431365
transform -1 0 162064 0 -1 4704
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _226_
timestamp 1698431365
transform 1 0 162512 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _227_
timestamp 1698431365
transform -1 0 165648 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _228_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 132720 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _229_
timestamp 1698431365
transform 1 0 134848 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _230_
timestamp 1698431365
transform 1 0 137200 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _231_
timestamp 1698431365
transform -1 0 96432 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _232_
timestamp 1698431365
transform -1 0 101024 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _233_
timestamp 1698431365
transform -1 0 104720 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _234_
timestamp 1698431365
transform -1 0 109200 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _235_
timestamp 1698431365
transform -1 0 112672 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _236_
timestamp 1698431365
transform -1 0 117040 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _237_
timestamp 1698431365
transform 1 0 117824 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _238_
timestamp 1698431365
transform -1 0 124656 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _239_
timestamp 1698431365
transform -1 0 129248 0 1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _240_
timestamp 1698431365
transform 1 0 131712 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _241_
timestamp 1698431365
transform 1 0 134960 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _242_
timestamp 1698431365
transform -1 0 140672 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _243_
timestamp 1698431365
transform 1 0 138768 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _252_
timestamp 1698431365
transform -1 0 93520 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _253_
timestamp 1698431365
transform -1 0 98112 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _254_
timestamp 1698431365
transform -1 0 101808 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _255_
timestamp 1698431365
transform -1 0 106288 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _256_
timestamp 1698431365
transform -1 0 109872 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _257_
timestamp 1698431365
transform -1 0 114128 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _258_
timestamp 1698431365
transform -1 0 118272 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _259_
timestamp 1698431365
transform -1 0 121968 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _260_
timestamp 1698431365
transform -1 0 126336 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _261_
timestamp 1698431365
transform -1 0 6160 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _262_
timestamp 1698431365
transform 1 0 49952 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _263_
timestamp 1698431365
transform 1 0 52640 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _264_
timestamp 1698431365
transform 1 0 55328 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _265_
timestamp 1698431365
transform 1 0 58016 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _266_
timestamp 1698431365
transform 1 0 60704 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _267_
timestamp 1698431365
transform 1 0 63392 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _268_
timestamp 1698431365
transform 1 0 66080 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _269_
timestamp 1698431365
transform 1 0 68768 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__108__A4 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 164752 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__110__B2
timestamp 1698431365
transform 1 0 135072 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__111__I
timestamp 1698431365
transform 1 0 131264 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__112__B2
timestamp 1698431365
transform -1 0 149184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__112__C1
timestamp 1698431365
transform 1 0 147616 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__113__A4
timestamp 1698431365
transform -1 0 147392 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__115__A2
timestamp 1698431365
transform -1 0 166992 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__116__A4
timestamp 1698431365
transform 1 0 164416 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__118__B2
timestamp 1698431365
transform -1 0 136416 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__119__I
timestamp 1698431365
transform 1 0 130816 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__120__B2
timestamp 1698431365
transform -1 0 153440 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__120__C1
timestamp 1698431365
transform 1 0 153664 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__121__A4
timestamp 1698431365
transform 1 0 154000 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__123__A2
timestamp 1698431365
transform -1 0 165200 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__124__A4
timestamp 1698431365
transform 1 0 163296 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__126__B2
timestamp 1698431365
transform -1 0 137984 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__127__I
timestamp 1698431365
transform 1 0 132608 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__128__B2
timestamp 1698431365
transform -1 0 150192 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__128__C1
timestamp 1698431365
transform 1 0 150080 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__129__A4
timestamp 1698431365
transform 1 0 155008 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__131__A2
timestamp 1698431365
transform -1 0 164192 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__132__A4
timestamp 1698431365
transform 1 0 162960 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__134__B2
timestamp 1698431365
transform -1 0 138544 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__136__B2
timestamp 1698431365
transform -1 0 154896 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__136__C1
timestamp 1698431365
transform 1 0 155120 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__137__A4
timestamp 1698431365
transform 1 0 150752 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__138__A3
timestamp 1698431365
transform 1 0 159936 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__139__A2
timestamp 1698431365
transform -1 0 163856 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__139__B
timestamp 1698431365
transform 1 0 160608 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__140__A4
timestamp 1698431365
transform -1 0 161168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__142__A1
timestamp 1698431365
transform -1 0 134624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__142__A2
timestamp 1698431365
transform 1 0 138656 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__142__B2
timestamp 1698431365
transform -1 0 139216 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__144__A1
timestamp 1698431365
transform -1 0 135856 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__145__A1
timestamp 1698431365
transform 1 0 138096 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__146__I
timestamp 1698431365
transform 1 0 139776 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__147__I
timestamp 1698431365
transform 1 0 149184 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__149__I
timestamp 1698431365
transform -1 0 147616 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__151__I
timestamp 1698431365
transform 1 0 147840 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__154__I
timestamp 1698431365
transform 1 0 138208 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__159__I
timestamp 1698431365
transform 1 0 148176 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__162__I
timestamp 1698431365
transform 1 0 140336 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__163__A4
timestamp 1698431365
transform -1 0 147504 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__167__A1
timestamp 1698431365
transform 1 0 146832 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__167__A2
timestamp 1698431365
transform 1 0 146160 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__168__I
timestamp 1698431365
transform -1 0 158032 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__169__A2
timestamp 1698431365
transform 1 0 154224 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__172__I
timestamp 1698431365
transform 1 0 160832 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__173__A2
timestamp 1698431365
transform 1 0 154672 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__180__A4
timestamp 1698431365
transform 1 0 154000 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__181__A2
timestamp 1698431365
transform 1 0 147840 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__184__I
timestamp 1698431365
transform -1 0 133504 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__185__B2
timestamp 1698431365
transform -1 0 143136 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__185__C1
timestamp 1698431365
transform -1 0 142912 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__188__A4
timestamp 1698431365
transform 1 0 153776 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__192__A4
timestamp 1698431365
transform 1 0 157920 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__195__I
timestamp 1698431365
transform 1 0 133728 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__196__B2
timestamp 1698431365
transform 1 0 145376 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__196__C1
timestamp 1698431365
transform 1 0 145824 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__197__A4
timestamp 1698431365
transform 1 0 152768 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__200__A4
timestamp 1698431365
transform -1 0 157248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__203__I
timestamp 1698431365
transform 1 0 135296 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__204__B2
timestamp 1698431365
transform 1 0 144256 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__204__C1
timestamp 1698431365
transform 1 0 145824 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__206__A4
timestamp 1698431365
transform 1 0 156128 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__210__A2
timestamp 1698431365
transform 1 0 165536 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__212__A4
timestamp 1698431365
transform -1 0 157808 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__214__B2
timestamp 1698431365
transform 1 0 140560 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__215__I
timestamp 1698431365
transform 1 0 130032 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__216__I
timestamp 1698431365
transform 1 0 135520 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__B2
timestamp 1698431365
transform -1 0 148848 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__C1
timestamp 1698431365
transform -1 0 148400 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__223__A4
timestamp 1698431365
transform 1 0 150304 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__224__I
timestamp 1698431365
transform 1 0 161056 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__226__I
timestamp 1698431365
transform 1 0 162288 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__A2
timestamp 1698431365
transform 1 0 165648 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__228__CLK
timestamp 1698431365
transform 1 0 136192 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__228__D
timestamp 1698431365
transform -1 0 132720 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__229__CLK
timestamp 1698431365
transform 1 0 134400 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__229__D
timestamp 1698431365
transform 1 0 133952 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__230__CLK
timestamp 1698431365
transform 1 0 136752 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__230__D
timestamp 1698431365
transform 1 0 136304 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__231__CLK
timestamp 1698431365
transform 1 0 96656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__231__D
timestamp 1698431365
transform 1 0 97104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__232__CLK
timestamp 1698431365
transform 1 0 101248 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__232__D
timestamp 1698431365
transform 1 0 101696 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__233__CLK
timestamp 1698431365
transform 1 0 104944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__233__D
timestamp 1698431365
transform 1 0 105392 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__234__CLK
timestamp 1698431365
transform 1 0 109424 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__234__D
timestamp 1698431365
transform 1 0 109872 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__235__CLK
timestamp 1698431365
transform 1 0 113344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__235__D
timestamp 1698431365
transform 1 0 112896 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__236__CLK
timestamp 1698431365
transform 1 0 113568 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__236__D
timestamp 1698431365
transform 1 0 117264 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__237__CLK
timestamp 1698431365
transform 1 0 117600 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__237__D
timestamp 1698431365
transform 1 0 121296 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__238__CLK
timestamp 1698431365
transform 1 0 125328 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__238__D
timestamp 1698431365
transform 1 0 124880 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__239__CLK
timestamp 1698431365
transform 1 0 129920 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__239__D
timestamp 1698431365
transform 1 0 129472 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__240__CLK
timestamp 1698431365
transform -1 0 135296 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__241__CLK
timestamp 1698431365
transform 1 0 135072 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__242__CLK
timestamp 1698431365
transform 1 0 137200 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__243__CLK
timestamp 1698431365
transform -1 0 138768 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__252__I
timestamp 1698431365
transform 1 0 93744 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__253__I
timestamp 1698431365
transform 1 0 98336 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__254__I
timestamp 1698431365
transform 1 0 102032 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__255__I
timestamp 1698431365
transform 1 0 106512 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__256__I
timestamp 1698431365
transform 1 0 110768 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__257__I
timestamp 1698431365
transform 1 0 114352 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__258__I
timestamp 1698431365
transform 1 0 118496 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__259__I
timestamp 1698431365
transform 1 0 122192 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__260__I
timestamp 1698431365
transform 1 0 126560 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__261__I
timestamp 1698431365
transform 1 0 6384 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__262__I
timestamp 1698431365
transform 1 0 49728 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__263__I
timestamp 1698431365
transform 1 0 52080 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__264__I
timestamp 1698431365
transform 1 0 55104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__265__I
timestamp 1698431365
transform 1 0 57792 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__266__I
timestamp 1698431365
transform 1 0 59920 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__267__I
timestamp 1698431365
transform 1 0 63168 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__268__I
timestamp 1698431365
transform 1 0 65856 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__269__I
timestamp 1698431365
transform 1 0 68544 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 118720 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_1_0__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 117152 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_1_1__f_wb_clk_i_I
timestamp 1698431365
transform 1 0 130480 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform -1 0 89712 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 92736 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform -1 0 95088 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform -1 0 97776 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform -1 0 100352 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform -1 0 103152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform -1 0 105840 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform -1 0 107968 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform -1 0 111776 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform -1 0 113904 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform -1 0 116592 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform -1 0 119392 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698431365
transform -1 0 121968 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698431365
transform -1 0 124656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698431365
transform -1 0 127008 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698431365
transform -1 0 130032 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698431365
transform -1 0 132720 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1698431365
transform -1 0 135408 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1698431365
transform -1 0 138432 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1698431365
transform -1 0 140784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1698431365
transform -1 0 143472 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1698431365
transform -1 0 146048 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1698431365
transform -1 0 147952 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1698431365
transform 1 0 155680 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1698431365
transform 1 0 156576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1698431365
transform -1 0 157472 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1698431365
transform -1 0 159600 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1698431365
transform -1 0 162064 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1698431365
transform -1 0 165088 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1698431365
transform -1 0 167664 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1698431365
transform -1 0 170352 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1698431365
transform -1 0 172704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1698431365
transform -1 0 175728 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input34_I
timestamp 1698431365
transform -1 0 178416 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input35_I
timestamp 1698431365
transform -1 0 181104 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input36_I
timestamp 1698431365
transform -1 0 184128 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input37_I
timestamp 1698431365
transform -1 0 186480 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input38_I
timestamp 1698431365
transform -1 0 189168 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input39_I
timestamp 1698431365
transform -1 0 191744 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input40_I
timestamp 1698431365
transform -1 0 194544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input41_I
timestamp 1698431365
transform -1 0 197232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input42_I
timestamp 1698431365
transform -1 0 199360 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input43_I
timestamp 1698431365
transform -1 0 203168 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input44_I
timestamp 1698431365
transform -1 0 205296 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input45_I
timestamp 1698431365
transform -1 0 207984 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input46_I
timestamp 1698431365
transform -1 0 210784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input47_I
timestamp 1698431365
transform -1 0 213360 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input48_I
timestamp 1698431365
transform -1 0 216048 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input49_I
timestamp 1698431365
transform -1 0 156240 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input50_I
timestamp 1698431365
transform -1 0 160272 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input51_I
timestamp 1698431365
transform -1 0 164304 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input52_I
timestamp 1698431365
transform 1 0 168672 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input53_I
timestamp 1698431365
transform 1 0 172480 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input54_I
timestamp 1698431365
transform 1 0 176288 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input55_I
timestamp 1698431365
transform -1 0 180320 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input56_I
timestamp 1698431365
transform -1 0 184128 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input57_I
timestamp 1698431365
transform -1 0 187936 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input58_I
timestamp 1698431365
transform -1 0 192528 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input59_I
timestamp 1698431365
transform -1 0 196560 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input60_I
timestamp 1698431365
transform -1 0 200592 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input61_I
timestamp 1698431365
transform -1 0 204624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input62_I
timestamp 1698431365
transform -1 0 208656 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input63_I
timestamp 1698431365
transform -1 0 212688 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input64_I
timestamp 1698431365
transform -1 0 216720 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input65_I
timestamp 1698431365
transform -1 0 11088 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input66_I
timestamp 1698431365
transform -1 0 15120 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input67_I
timestamp 1698431365
transform -1 0 19152 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input68_I
timestamp 1698431365
transform -1 0 23184 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input69_I
timestamp 1698431365
transform 1 0 27776 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input70_I
timestamp 1698431365
transform 1 0 31584 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input71_I
timestamp 1698431365
transform 1 0 35392 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input72_I
timestamp 1698431365
transform 1 0 39200 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input73_I
timestamp 1698431365
transform -1 0 43232 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input74_I
timestamp 1698431365
transform -1 0 79632 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input75_I
timestamp 1698431365
transform -1 0 83664 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input76_I
timestamp 1698431365
transform -1 0 123984 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input77_I
timestamp 1698431365
transform -1 0 128016 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input78_I
timestamp 1698431365
transform -1 0 132048 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input79_I
timestamp 1698431365
transform -1 0 136080 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input80_I
timestamp 1698431365
transform -1 0 140112 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input81_I
timestamp 1698431365
transform -1 0 144144 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input82_I
timestamp 1698431365
transform -1 0 87696 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input83_I
timestamp 1698431365
transform -1 0 91728 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input84_I
timestamp 1698431365
transform -1 0 95760 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input85_I
timestamp 1698431365
transform 1 0 100128 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input86_I
timestamp 1698431365
transform 1 0 103936 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input87_I
timestamp 1698431365
transform 1 0 107744 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input88_I
timestamp 1698431365
transform -1 0 111776 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input89_I
timestamp 1698431365
transform -1 0 115584 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input90_I
timestamp 1698431365
transform -1 0 119392 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input91_I
timestamp 1698431365
transform -1 0 7056 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output92_I
timestamp 1698431365
transform -1 0 31584 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output93_I
timestamp 1698431365
transform 1 0 33152 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output94_I
timestamp 1698431365
transform 1 0 35616 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output95_I
timestamp 1698431365
transform -1 0 39312 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output96_I
timestamp 1698431365
transform -1 0 43008 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output97_I
timestamp 1698431365
transform 1 0 44464 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output98_I
timestamp 1698431365
transform 1 0 46928 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output99_I
timestamp 1698431365
transform -1 0 50624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output100_I
timestamp 1698431365
transform 1 0 52528 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output110_I
timestamp 1698431365
transform -1 0 77280 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output111_I
timestamp 1698431365
transform -1 0 79632 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output112_I
timestamp 1698431365
transform 1 0 81312 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output113_I
timestamp 1698431365
transform -1 0 85008 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output114_I
timestamp 1698431365
transform 1 0 88032 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output115_I
timestamp 1698431365
transform 1 0 88928 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output116_I
timestamp 1698431365
transform 1 0 153216 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output117_I
timestamp 1698431365
transform -1 0 152208 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output118_I
timestamp 1698431365
transform 1 0 50512 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output119_I
timestamp 1698431365
transform 1 0 55104 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output120_I
timestamp 1698431365
transform 1 0 58912 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output121_I
timestamp 1698431365
transform 1 0 62720 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output122_I
timestamp 1698431365
transform 1 0 66528 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output123_I
timestamp 1698431365
transform 1 0 70336 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output124_I
timestamp 1698431365
transform 1 0 74144 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output125_I
timestamp 1698431365
transform -1 0 78960 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 119168 0 -1 37632
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_wb_clk_i
timestamp 1698431365
transform -1 0 116928 0 -1 32928
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_wb_clk_i
timestamp 1698431365
transform 1 0 130928 0 1 36064
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_36 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_44 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6272 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_49 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6832 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_65 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 8624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_67
timestamp 1698431365
transform 1 0 8848 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_74
timestamp 1698431365
transform 1 0 9632 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_90
timestamp 1698431365
transform 1 0 11424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_92
timestamp 1698431365
transform 1 0 11648 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_97 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12208 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_101
timestamp 1698431365
transform 1 0 12656 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_104
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_112
timestamp 1698431365
transform 1 0 13888 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_116
timestamp 1698431365
transform 1 0 14336 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_121
timestamp 1698431365
transform 1 0 14896 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_129
timestamp 1698431365
transform 1 0 15792 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_133
timestamp 1698431365
transform 1 0 16240 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_135
timestamp 1698431365
transform 1 0 16464 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_138
timestamp 1698431365
transform 1 0 16800 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_140
timestamp 1698431365
transform 1 0 17024 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_145
timestamp 1698431365
transform 1 0 17584 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_161
timestamp 1698431365
transform 1 0 19376 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_169
timestamp 1698431365
transform 1 0 20272 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_172
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_188
timestamp 1698431365
transform 1 0 22400 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_193
timestamp 1698431365
transform 1 0 22960 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_201
timestamp 1698431365
transform 1 0 23856 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_203
timestamp 1698431365
transform 1 0 24080 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_206
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_210
timestamp 1698431365
transform 1 0 24864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_212
timestamp 1698431365
transform 1 0 25088 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_217
timestamp 1698431365
transform 1 0 25648 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_233
timestamp 1698431365
transform 1 0 27440 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_237
timestamp 1698431365
transform 1 0 27888 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_266
timestamp 1698431365
transform 1 0 31136 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_270
timestamp 1698431365
transform 1 0 31584 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_274
timestamp 1698431365
transform 1 0 32032 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_278
timestamp 1698431365
transform 1 0 32480 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_308
timestamp 1698431365
transform 1 0 35840 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_335
timestamp 1698431365
transform 1 0 38864 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_339
timestamp 1698431365
transform 1 0 39312 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_368
timestamp 1698431365
transform 1 0 42560 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_372
timestamp 1698431365
transform 1 0 43008 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_376
timestamp 1698431365
transform 1 0 43456 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_380
timestamp 1698431365
transform 1 0 43904 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_407
timestamp 1698431365
transform 1 0 46928 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_436
timestamp 1698431365
transform 1 0 50176 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_440
timestamp 1698431365
transform 1 0 50624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_444
timestamp 1698431365
transform 1 0 51072 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_448
timestamp 1698431365
transform 1 0 51520 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_504
timestamp 1698431365
transform 1 0 57792 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_508
timestamp 1698431365
transform 1 0 58240 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_512
timestamp 1698431365
transform 1 0 58688 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_516
timestamp 1698431365
transform 1 0 59136 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_546
timestamp 1698431365
transform 1 0 62496 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_548
timestamp 1698431365
transform 1 0 62720 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_575
timestamp 1698431365
transform 1 0 65744 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_577
timestamp 1698431365
transform 1 0 65968 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_606
timestamp 1698431365
transform 1 0 69216 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_610
timestamp 1698431365
transform 1 0 69664 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_614
timestamp 1698431365
transform 1 0 70112 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_618
timestamp 1698431365
transform 1 0 70560 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_674
timestamp 1698431365
transform 1 0 76832 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_678
timestamp 1698431365
transform 1 0 77280 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_682
timestamp 1698431365
transform 1 0 77728 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_686
timestamp 1698431365
transform 1 0 78176 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_716
timestamp 1698431365
transform 1 0 81536 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_743
timestamp 1698431365
transform 1 0 84560 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_747
timestamp 1698431365
transform 1 0 85008 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_750
timestamp 1698431365
transform 1 0 85344 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_754
timestamp 1698431365
transform 1 0 85792 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_784
timestamp 1698431365
transform 1 0 89152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_786
timestamp 1698431365
transform 1 0 89376 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_795
timestamp 1698431365
transform 1 0 90384 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_811
timestamp 1698431365
transform 1 0 92176 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_813
timestamp 1698431365
transform 1 0 92400 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_824
timestamp 1698431365
transform 1 0 93632 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_832
timestamp 1698431365
transform 1 0 94528 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_834
timestamp 1698431365
transform 1 0 94752 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_843
timestamp 1698431365
transform 1 0 95760 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_847
timestamp 1698431365
transform 1 0 96208 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_849
timestamp 1698431365
transform 1 0 96432 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_852
timestamp 1698431365
transform 1 0 96768 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_856
timestamp 1698431365
transform 1 0 97216 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_858
timestamp 1698431365
transform 1 0 97440 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_867
timestamp 1698431365
transform 1 0 98448 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_875
timestamp 1698431365
transform 1 0 99344 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_879
timestamp 1698431365
transform 1 0 99792 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_881
timestamp 1698431365
transform 1 0 100016 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_892
timestamp 1698431365
transform 1 0 101248 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_900
timestamp 1698431365
transform 1 0 102144 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_904
timestamp 1698431365
transform 1 0 102592 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_906
timestamp 1698431365
transform 1 0 102816 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_915
timestamp 1698431365
transform 1 0 103824 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_917
timestamp 1698431365
transform 1 0 104048 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_920
timestamp 1698431365
transform 1 0 104384 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_928
timestamp 1698431365
transform 1 0 105280 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_930
timestamp 1698431365
transform 1 0 105504 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_939
timestamp 1698431365
transform 1 0 106512 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_947
timestamp 1698431365
transform 1 0 107408 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_949
timestamp 1698431365
transform 1 0 107632 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_954
timestamp 1698431365
transform 1 0 108192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_956
timestamp 1698431365
transform 1 0 108416 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_963
timestamp 1698431365
transform 1 0 109200 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_979
timestamp 1698431365
transform 1 0 110992 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_983
timestamp 1698431365
transform 1 0 111440 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_994
timestamp 1698431365
transform 1 0 112672 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1002
timestamp 1698431365
transform 1 0 113568 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_1011
timestamp 1698431365
transform 1 0 114576 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1019
timestamp 1698431365
transform 1 0 115472 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_1022
timestamp 1698431365
transform 1 0 115808 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1026
timestamp 1698431365
transform 1 0 116256 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_1035
timestamp 1698431365
transform 1 0 117264 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1051
timestamp 1698431365
transform 1 0 119056 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_1062
timestamp 1698431365
transform 1 0 120288 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_1070
timestamp 1698431365
transform 1 0 121184 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1074
timestamp 1698431365
transform 1 0 121632 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_1083
timestamp 1698431365
transform 1 0 122640 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1087
timestamp 1698431365
transform 1 0 123088 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_1090
timestamp 1698431365
transform 1 0 123424 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1098
timestamp 1698431365
transform 1 0 124320 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_1107
timestamp 1698431365
transform 1 0 125328 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_1115
timestamp 1698431365
transform 1 0 126224 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1119
timestamp 1698431365
transform 1 0 126672 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1124
timestamp 1698431365
transform 1 0 127232 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_1131
timestamp 1698431365
transform 1 0 128016 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1155
timestamp 1698431365
transform 1 0 130704 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_1158
timestamp 1698431365
transform 1 0 131040 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_1166
timestamp 1698431365
transform 1 0 131936 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1170
timestamp 1698431365
transform 1 0 132384 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_1179
timestamp 1698431365
transform 1 0 133392 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1187
timestamp 1698431365
transform 1 0 134288 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1189
timestamp 1698431365
transform 1 0 134512 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1192
timestamp 1698431365
transform 1 0 134848 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1194
timestamp 1698431365
transform 1 0 135072 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_1203
timestamp 1698431365
transform 1 0 136080 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1219
timestamp 1698431365
transform 1 0 137872 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1221
timestamp 1698431365
transform 1 0 138096 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_1232
timestamp 1698431365
transform 1 0 139328 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1240
timestamp 1698431365
transform 1 0 140224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1242
timestamp 1698431365
transform 1 0 140448 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_1251
timestamp 1698431365
transform 1 0 141456 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1255
timestamp 1698431365
transform 1 0 141904 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1257
timestamp 1698431365
transform 1 0 142128 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1260
timestamp 1698431365
transform 1 0 142464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1264
timestamp 1698431365
transform 1 0 142912 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1266
timestamp 1698431365
transform 1 0 143136 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_1275
timestamp 1698431365
transform 1 0 144144 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_1283
timestamp 1698431365
transform 1 0 145040 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1287
timestamp 1698431365
transform 1 0 145488 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1289
timestamp 1698431365
transform 1 0 145712 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1300
timestamp 1698431365
transform 1 0 146944 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1302
timestamp 1698431365
transform 1 0 147168 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1305
timestamp 1698431365
transform 1 0 147504 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1309
timestamp 1698431365
transform 1 0 147952 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1313
timestamp 1698431365
transform 1 0 148400 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1323
timestamp 1698431365
transform 1 0 149520 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1325
timestamp 1698431365
transform 1 0 149744 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1328
timestamp 1698431365
transform 1 0 150080 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1332
timestamp 1698431365
transform 1 0 150528 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1341
timestamp 1698431365
transform 1 0 151536 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1343
timestamp 1698431365
transform 1 0 151760 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1359
timestamp 1698431365
transform 1 0 153552 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1376
timestamp 1698431365
transform 1 0 155456 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1380
timestamp 1698431365
transform 1 0 155904 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1384
timestamp 1698431365
transform 1 0 156352 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_1388
timestamp 1698431365
transform 1 0 156800 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_1402
timestamp 1698431365
transform 1 0 158368 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1410
timestamp 1698431365
transform 1 0 159264 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_1419
timestamp 1698431365
transform 1 0 160272 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1427
timestamp 1698431365
transform 1 0 161168 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1430
timestamp 1698431365
transform 1 0 161504 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1432
timestamp 1698431365
transform 1 0 161728 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1435
timestamp 1698431365
transform 1 0 162064 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_1451
timestamp 1698431365
transform 1 0 163856 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1459
timestamp 1698431365
transform 1 0 164752 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_1470
timestamp 1698431365
transform 1 0 165984 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_1478
timestamp 1698431365
transform 1 0 166880 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1482
timestamp 1698431365
transform 1 0 167328 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_1491
timestamp 1698431365
transform 1 0 168336 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1495
timestamp 1698431365
transform 1 0 168784 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_1498
timestamp 1698431365
transform 1 0 169120 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1506
timestamp 1698431365
transform 1 0 170016 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_1515
timestamp 1698431365
transform 1 0 171024 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_1523
timestamp 1698431365
transform 1 0 171920 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1527
timestamp 1698431365
transform 1 0 172368 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1532
timestamp 1698431365
transform 1 0 172928 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_1539
timestamp 1698431365
transform 1 0 173712 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1563
timestamp 1698431365
transform 1 0 176400 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_1566
timestamp 1698431365
transform 1 0 176736 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_1574
timestamp 1698431365
transform 1 0 177632 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1578
timestamp 1698431365
transform 1 0 178080 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_1587
timestamp 1698431365
transform 1 0 179088 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1595
timestamp 1698431365
transform 1 0 179984 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1597
timestamp 1698431365
transform 1 0 180208 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1600
timestamp 1698431365
transform 1 0 180544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1602
timestamp 1698431365
transform 1 0 180768 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_1611
timestamp 1698431365
transform 1 0 181776 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1627
timestamp 1698431365
transform 1 0 183568 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1629
timestamp 1698431365
transform 1 0 183792 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_1640
timestamp 1698431365
transform 1 0 185024 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1648
timestamp 1698431365
transform 1 0 185920 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1650
timestamp 1698431365
transform 1 0 186144 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_1659
timestamp 1698431365
transform 1 0 187152 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1663
timestamp 1698431365
transform 1 0 187600 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1665
timestamp 1698431365
transform 1 0 187824 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_1668
timestamp 1698431365
transform 1 0 188160 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1672
timestamp 1698431365
transform 1 0 188608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1674
timestamp 1698431365
transform 1 0 188832 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_1683
timestamp 1698431365
transform 1 0 189840 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_1691
timestamp 1698431365
transform 1 0 190736 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1695
timestamp 1698431365
transform 1 0 191184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1697
timestamp 1698431365
transform 1 0 191408 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_1708
timestamp 1698431365
transform 1 0 192640 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_1716
timestamp 1698431365
transform 1 0 193536 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1720
timestamp 1698431365
transform 1 0 193984 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1722
timestamp 1698431365
transform 1 0 194208 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1731
timestamp 1698431365
transform 1 0 195216 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1733
timestamp 1698431365
transform 1 0 195440 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_1736
timestamp 1698431365
transform 1 0 195776 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1744
timestamp 1698431365
transform 1 0 196672 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1746
timestamp 1698431365
transform 1 0 196896 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_1757
timestamp 1698431365
transform 1 0 198128 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1765
timestamp 1698431365
transform 1 0 199024 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1770
timestamp 1698431365
transform 1 0 199584 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1772
timestamp 1698431365
transform 1 0 199808 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_1781
timestamp 1698431365
transform 1 0 200816 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1797
timestamp 1698431365
transform 1 0 202608 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1799
timestamp 1698431365
transform 1 0 202832 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_1812
timestamp 1698431365
transform 1 0 204288 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1816
timestamp 1698431365
transform 1 0 204736 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1818
timestamp 1698431365
transform 1 0 204960 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_1829
timestamp 1698431365
transform 1 0 206192 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1833
timestamp 1698431365
transform 1 0 206640 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1835
timestamp 1698431365
transform 1 0 206864 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_1838
timestamp 1698431365
transform 1 0 207200 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1842
timestamp 1698431365
transform 1 0 207648 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_1853
timestamp 1698431365
transform 1 0 208880 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_1861
timestamp 1698431365
transform 1 0 209776 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1865
timestamp 1698431365
transform 1 0 210224 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1867
timestamp 1698431365
transform 1 0 210448 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_1880
timestamp 1698431365
transform 1 0 211904 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1888
timestamp 1698431365
transform 1 0 212800 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1890
timestamp 1698431365
transform 1 0 213024 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_1901
timestamp 1698431365
transform 1 0 214256 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1903
timestamp 1698431365
transform 1 0 214480 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_1906
timestamp 1698431365
transform 1 0 214816 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1914
timestamp 1698431365
transform 1 0 215712 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_1925
timestamp 1698431365
transform 1 0 216944 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_1933
timestamp 1698431365
transform 1 0 217840 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_1937
timestamp 1698431365
transform 1 0 218288 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_2
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_18
timestamp 1698431365
transform 1 0 3360 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_20
timestamp 1698431365
transform 1 0 3584 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_47
timestamp 1698431365
transform 1 0 6608 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_63
timestamp 1698431365
transform 1 0 8400 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_67
timestamp 1698431365
transform 1 0 8848 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_69
timestamp 1698431365
transform 1 0 9072 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698431365
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_142
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_206
timestamp 1698431365
transform 1 0 24416 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_212
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_244
timestamp 1698431365
transform 1 0 28672 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_252
timestamp 1698431365
transform 1 0 29568 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_282
timestamp 1698431365
transform 1 0 32928 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_286
timestamp 1698431365
transform 1 0 33376 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_302
timestamp 1698431365
transform 1 0 35168 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_308
timestamp 1698431365
transform 1 0 35840 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_340
timestamp 1698431365
transform 1 0 39424 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_348
timestamp 1698431365
transform 1 0 40320 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_352
timestamp 1698431365
transform 1 0 40768 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_356
timestamp 1698431365
transform 1 0 41216 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_383
timestamp 1698431365
transform 1 0 44240 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_387
timestamp 1698431365
transform 1 0 44688 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_403
timestamp 1698431365
transform 1 0 46480 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_409
timestamp 1698431365
transform 1 0 47152 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_417
timestamp 1698431365
transform 1 0 48048 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_419
timestamp 1698431365
transform 1 0 48272 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_422
timestamp 1698431365
transform 1 0 48608 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_426
timestamp 1698431365
transform 1 0 49056 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_428
timestamp 1698431365
transform 1 0 49280 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_455
timestamp 1698431365
transform 1 0 52304 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_459
timestamp 1698431365
transform 1 0 52752 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_475
timestamp 1698431365
transform 1 0 54544 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_483
timestamp 1698431365
transform 1 0 55440 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_487
timestamp 1698431365
transform 1 0 55888 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_489
timestamp 1698431365
transform 1 0 56112 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_492
timestamp 1698431365
transform 1 0 56448 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_500
timestamp 1698431365
transform 1 0 57344 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_527
timestamp 1698431365
transform 1 0 60368 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_559
timestamp 1698431365
transform 1 0 63952 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_562
timestamp 1698431365
transform 1 0 64288 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_594
timestamp 1698431365
transform 1 0 67872 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_596
timestamp 1698431365
transform 1 0 68096 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_623
timestamp 1698431365
transform 1 0 71120 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_627
timestamp 1698431365
transform 1 0 71568 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_629
timestamp 1698431365
transform 1 0 71792 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_632
timestamp 1698431365
transform 1 0 72128 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_664
timestamp 1698431365
transform 1 0 75712 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_668
timestamp 1698431365
transform 1 0 76160 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_695
timestamp 1698431365
transform 1 0 79184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_699
timestamp 1698431365
transform 1 0 79632 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_702
timestamp 1698431365
transform 1 0 79968 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_710
timestamp 1698431365
transform 1 0 80864 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_716
timestamp 1698431365
transform 1 0 81536 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_732
timestamp 1698431365
transform 1 0 83328 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_740
timestamp 1698431365
transform 1 0 84224 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_767
timestamp 1698431365
transform 1 0 87248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_769
timestamp 1698431365
transform 1 0 87472 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_772
timestamp 1698431365
transform 1 0 87808 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_776
timestamp 1698431365
transform 1 0 88256 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_780
timestamp 1698431365
transform 1 0 88704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_784
timestamp 1698431365
transform 1 0 89152 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_816
timestamp 1698431365
transform 1 0 92736 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_832
timestamp 1698431365
transform 1 0 94528 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_842
timestamp 1698431365
transform 1 0 95648 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_906
timestamp 1698431365
transform 1 0 102816 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_912
timestamp 1698431365
transform 1 0 103488 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_976
timestamp 1698431365
transform 1 0 110656 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_982
timestamp 1698431365
transform 1 0 111328 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_1046
timestamp 1698431365
transform 1 0 118496 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_1052
timestamp 1698431365
transform 1 0 119168 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_1116
timestamp 1698431365
transform 1 0 126336 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_1122
timestamp 1698431365
transform 1 0 127008 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_1154
timestamp 1698431365
transform 1 0 130592 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_1158
timestamp 1698431365
transform 1 0 131040 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_1162
timestamp 1698431365
transform 1 0 131488 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_1178
timestamp 1698431365
transform 1 0 133280 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_1184
timestamp 1698431365
transform 1 0 133952 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_1188
timestamp 1698431365
transform 1 0 134400 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_1192
timestamp 1698431365
transform 1 0 134848 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_1198
timestamp 1698431365
transform 1 0 135520 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_1206
timestamp 1698431365
transform 1 0 136416 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_1210
timestamp 1698431365
transform 1 0 136864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_1212
timestamp 1698431365
transform 1 0 137088 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_1262
timestamp 1698431365
transform 1 0 142688 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_1266
timestamp 1698431365
transform 1 0 143136 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_1370
timestamp 1698431365
transform 1 0 154784 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_1387
timestamp 1698431365
transform 1 0 156688 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_1395
timestamp 1698431365
transform 1 0 157584 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_1399
timestamp 1698431365
transform 1 0 158032 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_1402
timestamp 1698431365
transform 1 0 158368 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_1418
timestamp 1698431365
transform 1 0 160160 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_1422
timestamp 1698431365
transform 1 0 160608 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_1426
timestamp 1698431365
transform 1 0 161056 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_1435
timestamp 1698431365
transform 1 0 162064 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_1456
timestamp 1698431365
transform 1 0 164416 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_1464
timestamp 1698431365
transform 1 0 165312 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_1466
timestamp 1698431365
transform 1 0 165536 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_1469
timestamp 1698431365
transform 1 0 165872 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_1472
timestamp 1698431365
transform 1 0 166208 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_1536
timestamp 1698431365
transform 1 0 173376 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_1542
timestamp 1698431365
transform 1 0 174048 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_1606
timestamp 1698431365
transform 1 0 181216 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_1612
timestamp 1698431365
transform 1 0 181888 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_1676
timestamp 1698431365
transform 1 0 189056 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_1682
timestamp 1698431365
transform 1 0 189728 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_1746
timestamp 1698431365
transform 1 0 196896 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_1752
timestamp 1698431365
transform 1 0 197568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_1816
timestamp 1698431365
transform 1 0 204736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_1822
timestamp 1698431365
transform 1 0 205408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_1886
timestamp 1698431365
transform 1 0 212576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_1892
timestamp 1698431365
transform 1 0 213248 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_1924
timestamp 1698431365
transform 1 0 216832 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_1932
timestamp 1698431365
transform 1 0 217728 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_1936
timestamp 1698431365
transform 1 0 218176 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_43
timestamp 1698431365
transform 1 0 6160 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_47
timestamp 1698431365
transform 1 0 6608 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_79
timestamp 1698431365
transform 1 0 10192 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_95
timestamp 1698431365
transform 1 0 11984 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_103
timestamp 1698431365
transform 1 0 12880 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698431365
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698431365
transform 1 0 28336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698431365
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698431365
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_317
timestamp 1698431365
transform 1 0 36848 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_381
timestamp 1698431365
transform 1 0 44016 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_387
timestamp 1698431365
transform 1 0 44688 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_419
timestamp 1698431365
transform 1 0 48272 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_427
timestamp 1698431365
transform 1 0 49168 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_431
timestamp 1698431365
transform 1 0 49616 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_440
timestamp 1698431365
transform 1 0 50624 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_448
timestamp 1698431365
transform 1 0 51520 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_452
timestamp 1698431365
transform 1 0 51968 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_457
timestamp 1698431365
transform 1 0 52528 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_464
timestamp 1698431365
transform 1 0 53312 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_488
timestamp 1698431365
transform 1 0 56000 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_512
timestamp 1698431365
transform 1 0 58688 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_520
timestamp 1698431365
transform 1 0 59584 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_522
timestamp 1698431365
transform 1 0 59808 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_527
timestamp 1698431365
transform 1 0 60368 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_529
timestamp 1698431365
transform 1 0 60592 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_536
timestamp 1698431365
transform 1 0 61376 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_560
timestamp 1698431365
transform 1 0 64064 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_584
timestamp 1698431365
transform 1 0 66752 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_592
timestamp 1698431365
transform 1 0 67648 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_594
timestamp 1698431365
transform 1 0 67872 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_597
timestamp 1698431365
transform 1 0 68208 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_599
timestamp 1698431365
transform 1 0 68432 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_608
timestamp 1698431365
transform 1 0 69440 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_640
timestamp 1698431365
transform 1 0 73024 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_656
timestamp 1698431365
transform 1 0 74816 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_664
timestamp 1698431365
transform 1 0 75712 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_667
timestamp 1698431365
transform 1 0 76048 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_731
timestamp 1698431365
transform 1 0 83216 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_737
timestamp 1698431365
transform 1 0 83888 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_801
timestamp 1698431365
transform 1 0 91056 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_807
timestamp 1698431365
transform 1 0 91728 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_823
timestamp 1698431365
transform 1 0 93520 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_827
timestamp 1698431365
transform 1 0 93968 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_843
timestamp 1698431365
transform 1 0 95760 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_851
timestamp 1698431365
transform 1 0 96656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_855
timestamp 1698431365
transform 1 0 97104 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_864
timestamp 1698431365
transform 1 0 98112 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_868
timestamp 1698431365
transform 1 0 98560 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_872
timestamp 1698431365
transform 1 0 99008 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_874
timestamp 1698431365
transform 1 0 99232 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_877
timestamp 1698431365
transform 1 0 99568 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_885
timestamp 1698431365
transform 1 0 100464 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_897
timestamp 1698431365
transform 1 0 101808 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_901
timestamp 1698431365
transform 1 0 102256 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_917
timestamp 1698431365
transform 1 0 104048 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_925
timestamp 1698431365
transform 1 0 104944 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_937
timestamp 1698431365
transform 1 0 106288 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_941
timestamp 1698431365
transform 1 0 106736 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_947
timestamp 1698431365
transform 1 0 107408 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_955
timestamp 1698431365
transform 1 0 108304 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_959
timestamp 1698431365
transform 1 0 108752 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_975
timestamp 1698431365
transform 1 0 110544 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_979
timestamp 1698431365
transform 1 0 110992 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_995
timestamp 1698431365
transform 1 0 112784 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_1007
timestamp 1698431365
transform 1 0 114128 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_1011
timestamp 1698431365
transform 1 0 114576 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_1017
timestamp 1698431365
transform 1 0 115248 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_1033
timestamp 1698431365
transform 1 0 117040 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_1035
timestamp 1698431365
transform 1 0 117264 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_1044
timestamp 1698431365
transform 1 0 118272 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_1048
timestamp 1698431365
transform 1 0 118720 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_1064
timestamp 1698431365
transform 1 0 120512 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_1068
timestamp 1698431365
transform 1 0 120960 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_1077
timestamp 1698431365
transform 1 0 121968 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_1081
timestamp 1698431365
transform 1 0 122416 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_1087
timestamp 1698431365
transform 1 0 123088 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_1103
timestamp 1698431365
transform 1 0 124880 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_1107
timestamp 1698431365
transform 1 0 125328 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_1116
timestamp 1698431365
transform 1 0 126336 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_1120
timestamp 1698431365
transform 1 0 126784 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_1136
timestamp 1698431365
transform 1 0 128576 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_1144
timestamp 1698431365
transform 1 0 129472 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_1148
timestamp 1698431365
transform 1 0 129920 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_1157
timestamp 1698431365
transform 1 0 130928 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_1170
timestamp 1698431365
transform 1 0 132384 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_1174
timestamp 1698431365
transform 1 0 132832 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_1202
timestamp 1698431365
transform 1 0 135968 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_1213
timestamp 1698431365
transform 1 0 137200 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_1223
timestamp 1698431365
transform 1 0 138320 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_1284
timestamp 1698431365
transform 1 0 145152 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_1288
timestamp 1698431365
transform 1 0 145600 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_1292
timestamp 1698431365
transform 1 0 146048 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_1294
timestamp 1698431365
transform 1 0 146272 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_1353
timestamp 1698431365
transform 1 0 152880 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_1403
timestamp 1698431365
transform 1 0 158480 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_1411
timestamp 1698431365
transform 1 0 159376 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_1415
timestamp 1698431365
transform 1 0 159824 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_1417
timestamp 1698431365
transform 1 0 160048 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_1445
timestamp 1698431365
transform 1 0 163184 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_1475
timestamp 1698431365
transform 1 0 166544 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_1479
timestamp 1698431365
transform 1 0 166992 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_1495
timestamp 1698431365
transform 1 0 168784 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_1503
timestamp 1698431365
transform 1 0 169680 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_1507
timestamp 1698431365
transform 1 0 170128 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_1571
timestamp 1698431365
transform 1 0 177296 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_1577
timestamp 1698431365
transform 1 0 177968 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_1641
timestamp 1698431365
transform 1 0 185136 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_1647
timestamp 1698431365
transform 1 0 185808 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_1711
timestamp 1698431365
transform 1 0 192976 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_1717
timestamp 1698431365
transform 1 0 193648 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_1781
timestamp 1698431365
transform 1 0 200816 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_1787
timestamp 1698431365
transform 1 0 201488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_1851
timestamp 1698431365
transform 1 0 208656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_1857
timestamp 1698431365
transform 1 0 209328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_1921
timestamp 1698431365
transform 1 0 216496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_1927
timestamp 1698431365
transform 1 0 217168 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_1935
timestamp 1698431365
transform 1 0 218064 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_1937
timestamp 1698431365
transform 1 0 218288 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698431365
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698431365
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698431365
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698431365
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698431365
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_346
timestamp 1698431365
transform 1 0 40096 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_352
timestamp 1698431365
transform 1 0 40768 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_416
timestamp 1698431365
transform 1 0 47936 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_422
timestamp 1698431365
transform 1 0 48608 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_486
timestamp 1698431365
transform 1 0 55776 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_492
timestamp 1698431365
transform 1 0 56448 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_556
timestamp 1698431365
transform 1 0 63616 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_562
timestamp 1698431365
transform 1 0 64288 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_626
timestamp 1698431365
transform 1 0 71456 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_632
timestamp 1698431365
transform 1 0 72128 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_696
timestamp 1698431365
transform 1 0 79296 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_702
timestamp 1698431365
transform 1 0 79968 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_766
timestamp 1698431365
transform 1 0 87136 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_772
timestamp 1698431365
transform 1 0 87808 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_836
timestamp 1698431365
transform 1 0 94976 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_842
timestamp 1698431365
transform 1 0 95648 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_906
timestamp 1698431365
transform 1 0 102816 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_912
timestamp 1698431365
transform 1 0 103488 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_976
timestamp 1698431365
transform 1 0 110656 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_982
timestamp 1698431365
transform 1 0 111328 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_1046
timestamp 1698431365
transform 1 0 118496 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_1052
timestamp 1698431365
transform 1 0 119168 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_1116
timestamp 1698431365
transform 1 0 126336 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_1122
timestamp 1698431365
transform 1 0 127008 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_1186
timestamp 1698431365
transform 1 0 134176 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_1192
timestamp 1698431365
transform 1 0 134848 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_1196
timestamp 1698431365
transform 1 0 135296 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_1241
timestamp 1698431365
transform 1 0 140336 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_1245
timestamp 1698431365
transform 1 0 140784 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_1256
timestamp 1698431365
transform 1 0 142016 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_1262
timestamp 1698431365
transform 1 0 142688 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_1266
timestamp 1698431365
transform 1 0 143136 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_1268
timestamp 1698431365
transform 1 0 143360 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_1316
timestamp 1698431365
transform 1 0 148736 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_1320
timestamp 1698431365
transform 1 0 149184 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_1332
timestamp 1698431365
transform 1 0 150528 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_1336
timestamp 1698431365
transform 1 0 150976 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_1395
timestamp 1698431365
transform 1 0 157584 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_1399
timestamp 1698431365
transform 1 0 158032 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_1402
timestamp 1698431365
transform 1 0 158368 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_1406
timestamp 1698431365
transform 1 0 158816 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_1408
timestamp 1698431365
transform 1 0 159040 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_1434
timestamp 1698431365
transform 1 0 161952 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_1436
timestamp 1698431365
transform 1 0 162176 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_1464
timestamp 1698431365
transform 1 0 165312 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_1468
timestamp 1698431365
transform 1 0 165760 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_1472
timestamp 1698431365
transform 1 0 166208 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_1536
timestamp 1698431365
transform 1 0 173376 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_1542
timestamp 1698431365
transform 1 0 174048 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_1606
timestamp 1698431365
transform 1 0 181216 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_1612
timestamp 1698431365
transform 1 0 181888 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_1676
timestamp 1698431365
transform 1 0 189056 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_1682
timestamp 1698431365
transform 1 0 189728 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_1746
timestamp 1698431365
transform 1 0 196896 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_1752
timestamp 1698431365
transform 1 0 197568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_1816
timestamp 1698431365
transform 1 0 204736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_1822
timestamp 1698431365
transform 1 0 205408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_1886
timestamp 1698431365
transform 1 0 212576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_1892
timestamp 1698431365
transform 1 0 213248 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_1924
timestamp 1698431365
transform 1 0 216832 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_1932
timestamp 1698431365
transform 1 0 217728 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_1936
timestamp 1698431365
transform 1 0 218176 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698431365
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698431365
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698431365
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698431365
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_317
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_381
timestamp 1698431365
transform 1 0 44016 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_387
timestamp 1698431365
transform 1 0 44688 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_451
timestamp 1698431365
transform 1 0 51856 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_457
timestamp 1698431365
transform 1 0 52528 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_521
timestamp 1698431365
transform 1 0 59696 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_527
timestamp 1698431365
transform 1 0 60368 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_591
timestamp 1698431365
transform 1 0 67536 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_597
timestamp 1698431365
transform 1 0 68208 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_661
timestamp 1698431365
transform 1 0 75376 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_667
timestamp 1698431365
transform 1 0 76048 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_731
timestamp 1698431365
transform 1 0 83216 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_737
timestamp 1698431365
transform 1 0 83888 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_801
timestamp 1698431365
transform 1 0 91056 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_807
timestamp 1698431365
transform 1 0 91728 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_871
timestamp 1698431365
transform 1 0 98896 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_877
timestamp 1698431365
transform 1 0 99568 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_941
timestamp 1698431365
transform 1 0 106736 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_947
timestamp 1698431365
transform 1 0 107408 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_1011
timestamp 1698431365
transform 1 0 114576 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_1017
timestamp 1698431365
transform 1 0 115248 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_1081
timestamp 1698431365
transform 1 0 122416 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_1087
timestamp 1698431365
transform 1 0 123088 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_1151
timestamp 1698431365
transform 1 0 130256 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_1157
timestamp 1698431365
transform 1 0 130928 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_1165
timestamp 1698431365
transform 1 0 131824 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_1169
timestamp 1698431365
transform 1 0 132272 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_1216
timestamp 1698431365
transform 1 0 137536 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_1220
timestamp 1698431365
transform 1 0 137984 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_1224
timestamp 1698431365
transform 1 0 138432 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_1274
timestamp 1698431365
transform 1 0 144032 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_1288
timestamp 1698431365
transform 1 0 145600 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_1292
timestamp 1698431365
transform 1 0 146048 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_1294
timestamp 1698431365
transform 1 0 146272 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_1297
timestamp 1698431365
transform 1 0 146608 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_1301
timestamp 1698431365
transform 1 0 147056 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_1304
timestamp 1698431365
transform 1 0 147392 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_1361
timestamp 1698431365
transform 1 0 153776 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_1367
timestamp 1698431365
transform 1 0 154448 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_1394
timestamp 1698431365
transform 1 0 157472 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_1410
timestamp 1698431365
transform 1 0 159264 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_1414
timestamp 1698431365
transform 1 0 159712 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_1433
timestamp 1698431365
transform 1 0 161840 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_1437
timestamp 1698431365
transform 1 0 162288 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_1447
timestamp 1698431365
transform 1 0 163408 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_1459
timestamp 1698431365
transform 1 0 164752 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_1463
timestamp 1698431365
transform 1 0 165200 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_1495
timestamp 1698431365
transform 1 0 168784 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_1503
timestamp 1698431365
transform 1 0 169680 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_1507
timestamp 1698431365
transform 1 0 170128 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_1571
timestamp 1698431365
transform 1 0 177296 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_1577
timestamp 1698431365
transform 1 0 177968 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_1641
timestamp 1698431365
transform 1 0 185136 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_1647
timestamp 1698431365
transform 1 0 185808 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_1711
timestamp 1698431365
transform 1 0 192976 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_1717
timestamp 1698431365
transform 1 0 193648 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_1781
timestamp 1698431365
transform 1 0 200816 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_1787
timestamp 1698431365
transform 1 0 201488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_1851
timestamp 1698431365
transform 1 0 208656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_1857
timestamp 1698431365
transform 1 0 209328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_1921
timestamp 1698431365
transform 1 0 216496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_1927
timestamp 1698431365
transform 1 0 217168 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_1935
timestamp 1698431365
transform 1 0 218064 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_1937
timestamp 1698431365
transform 1 0 218288 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698431365
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698431365
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698431365
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698431365
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_346
timestamp 1698431365
transform 1 0 40096 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_352
timestamp 1698431365
transform 1 0 40768 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_416
timestamp 1698431365
transform 1 0 47936 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_422
timestamp 1698431365
transform 1 0 48608 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_486
timestamp 1698431365
transform 1 0 55776 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_492
timestamp 1698431365
transform 1 0 56448 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_556
timestamp 1698431365
transform 1 0 63616 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_562
timestamp 1698431365
transform 1 0 64288 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_626
timestamp 1698431365
transform 1 0 71456 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_632
timestamp 1698431365
transform 1 0 72128 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_696
timestamp 1698431365
transform 1 0 79296 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_702
timestamp 1698431365
transform 1 0 79968 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_766
timestamp 1698431365
transform 1 0 87136 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_772
timestamp 1698431365
transform 1 0 87808 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_836
timestamp 1698431365
transform 1 0 94976 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_842
timestamp 1698431365
transform 1 0 95648 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_906
timestamp 1698431365
transform 1 0 102816 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_912
timestamp 1698431365
transform 1 0 103488 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_976
timestamp 1698431365
transform 1 0 110656 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_982
timestamp 1698431365
transform 1 0 111328 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_1046
timestamp 1698431365
transform 1 0 118496 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_1052
timestamp 1698431365
transform 1 0 119168 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_1116
timestamp 1698431365
transform 1 0 126336 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_1122
timestamp 1698431365
transform 1 0 127008 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_1154
timestamp 1698431365
transform 1 0 130592 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_1256
timestamp 1698431365
transform 1 0 142016 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_1276
timestamp 1698431365
transform 1 0 144256 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_1325
timestamp 1698431365
transform 1 0 149744 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_1329
timestamp 1698431365
transform 1 0 150192 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_1359
timestamp 1698431365
transform 1 0 153552 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_1363
timestamp 1698431365
transform 1 0 154000 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_1367
timestamp 1698431365
transform 1 0 154448 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_1371
timestamp 1698431365
transform 1 0 154896 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_1375
timestamp 1698431365
transform 1 0 155344 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_1391
timestamp 1698431365
transform 1 0 157136 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_1399
timestamp 1698431365
transform 1 0 158032 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_1402
timestamp 1698431365
transform 1 0 158368 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_1418
timestamp 1698431365
transform 1 0 160160 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_1424
timestamp 1698431365
transform 1 0 160832 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_1434
timestamp 1698431365
transform 1 0 161952 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_1450
timestamp 1698431365
transform 1 0 163744 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_1454
timestamp 1698431365
transform 1 0 164192 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_1472
timestamp 1698431365
transform 1 0 166208 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_1536
timestamp 1698431365
transform 1 0 173376 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_1542
timestamp 1698431365
transform 1 0 174048 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_1606
timestamp 1698431365
transform 1 0 181216 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_1612
timestamp 1698431365
transform 1 0 181888 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_1676
timestamp 1698431365
transform 1 0 189056 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_1682
timestamp 1698431365
transform 1 0 189728 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_1746
timestamp 1698431365
transform 1 0 196896 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_1752
timestamp 1698431365
transform 1 0 197568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_1816
timestamp 1698431365
transform 1 0 204736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_1822
timestamp 1698431365
transform 1 0 205408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_1886
timestamp 1698431365
transform 1 0 212576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_1892
timestamp 1698431365
transform 1 0 213248 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_1924
timestamp 1698431365
transform 1 0 216832 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_1932
timestamp 1698431365
transform 1 0 217728 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_1936
timestamp 1698431365
transform 1 0 218176 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698431365
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698431365
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698431365
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698431365
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_317
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_381
timestamp 1698431365
transform 1 0 44016 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_387
timestamp 1698431365
transform 1 0 44688 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_451
timestamp 1698431365
transform 1 0 51856 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_457
timestamp 1698431365
transform 1 0 52528 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_521
timestamp 1698431365
transform 1 0 59696 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_527
timestamp 1698431365
transform 1 0 60368 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_591
timestamp 1698431365
transform 1 0 67536 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_597
timestamp 1698431365
transform 1 0 68208 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_661
timestamp 1698431365
transform 1 0 75376 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_667
timestamp 1698431365
transform 1 0 76048 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_731
timestamp 1698431365
transform 1 0 83216 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_737
timestamp 1698431365
transform 1 0 83888 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_801
timestamp 1698431365
transform 1 0 91056 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_807
timestamp 1698431365
transform 1 0 91728 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_871
timestamp 1698431365
transform 1 0 98896 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_877
timestamp 1698431365
transform 1 0 99568 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_941
timestamp 1698431365
transform 1 0 106736 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_947
timestamp 1698431365
transform 1 0 107408 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_1011
timestamp 1698431365
transform 1 0 114576 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_1017
timestamp 1698431365
transform 1 0 115248 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_1081
timestamp 1698431365
transform 1 0 122416 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_1087
timestamp 1698431365
transform 1 0 123088 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_1151
timestamp 1698431365
transform 1 0 130256 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_1157
timestamp 1698431365
transform 1 0 130928 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_1165
timestamp 1698431365
transform 1 0 131824 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_1169
timestamp 1698431365
transform 1 0 132272 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_1202
timestamp 1698431365
transform 1 0 135968 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_1206
timestamp 1698431365
transform 1 0 136416 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_1222
timestamp 1698431365
transform 1 0 138208 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_1259
timestamp 1698431365
transform 1 0 142352 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_1263
timestamp 1698431365
transform 1 0 142800 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_1265
timestamp 1698431365
transform 1 0 143024 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_1286
timestamp 1698431365
transform 1 0 145376 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_1294
timestamp 1698431365
transform 1 0 146272 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_1297
timestamp 1698431365
transform 1 0 146608 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_1305
timestamp 1698431365
transform 1 0 147504 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_1307
timestamp 1698431365
transform 1 0 147728 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_1350
timestamp 1698431365
transform 1 0 152544 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_1354
timestamp 1698431365
transform 1 0 152992 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_1358
timestamp 1698431365
transform 1 0 153440 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_1362
timestamp 1698431365
transform 1 0 153888 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_1364
timestamp 1698431365
transform 1 0 154112 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_1367
timestamp 1698431365
transform 1 0 154448 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_1371
timestamp 1698431365
transform 1 0 154896 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_1443
timestamp 1698431365
transform 1 0 162960 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_1475
timestamp 1698431365
transform 1 0 166544 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_1491
timestamp 1698431365
transform 1 0 168336 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_1499
timestamp 1698431365
transform 1 0 169232 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_1503
timestamp 1698431365
transform 1 0 169680 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_1507
timestamp 1698431365
transform 1 0 170128 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_1571
timestamp 1698431365
transform 1 0 177296 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_1577
timestamp 1698431365
transform 1 0 177968 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_1641
timestamp 1698431365
transform 1 0 185136 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_1647
timestamp 1698431365
transform 1 0 185808 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_1711
timestamp 1698431365
transform 1 0 192976 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_1717
timestamp 1698431365
transform 1 0 193648 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_1781
timestamp 1698431365
transform 1 0 200816 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_1787
timestamp 1698431365
transform 1 0 201488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_1851
timestamp 1698431365
transform 1 0 208656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_1857
timestamp 1698431365
transform 1 0 209328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_1921
timestamp 1698431365
transform 1 0 216496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_1927
timestamp 1698431365
transform 1 0 217168 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_1935
timestamp 1698431365
transform 1 0 218064 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_1937
timestamp 1698431365
transform 1 0 218288 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698431365
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698431365
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698431365
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698431365
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698431365
transform 1 0 32928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_346
timestamp 1698431365
transform 1 0 40096 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_352
timestamp 1698431365
transform 1 0 40768 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_416
timestamp 1698431365
transform 1 0 47936 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_422
timestamp 1698431365
transform 1 0 48608 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_486
timestamp 1698431365
transform 1 0 55776 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_492
timestamp 1698431365
transform 1 0 56448 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_556
timestamp 1698431365
transform 1 0 63616 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_562
timestamp 1698431365
transform 1 0 64288 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_626
timestamp 1698431365
transform 1 0 71456 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_632
timestamp 1698431365
transform 1 0 72128 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_696
timestamp 1698431365
transform 1 0 79296 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_702
timestamp 1698431365
transform 1 0 79968 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_766
timestamp 1698431365
transform 1 0 87136 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_772
timestamp 1698431365
transform 1 0 87808 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_836
timestamp 1698431365
transform 1 0 94976 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_842
timestamp 1698431365
transform 1 0 95648 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_906
timestamp 1698431365
transform 1 0 102816 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_912
timestamp 1698431365
transform 1 0 103488 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_976
timestamp 1698431365
transform 1 0 110656 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_982
timestamp 1698431365
transform 1 0 111328 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_1046
timestamp 1698431365
transform 1 0 118496 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_1052
timestamp 1698431365
transform 1 0 119168 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_1116
timestamp 1698431365
transform 1 0 126336 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_1122
timestamp 1698431365
transform 1 0 127008 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_1186
timestamp 1698431365
transform 1 0 134176 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_1224
timestamp 1698431365
transform 1 0 138432 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_1236
timestamp 1698431365
transform 1 0 139776 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_1238
timestamp 1698431365
transform 1 0 140000 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_1248
timestamp 1698431365
transform 1 0 141120 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_1256
timestamp 1698431365
transform 1 0 142016 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_1262
timestamp 1698431365
transform 1 0 142688 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_1294
timestamp 1698431365
transform 1 0 146272 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_1326
timestamp 1698431365
transform 1 0 149856 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_1364
timestamp 1698431365
transform 1 0 154112 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_1388
timestamp 1698431365
transform 1 0 156800 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_1392
timestamp 1698431365
transform 1 0 157248 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_1402
timestamp 1698431365
transform 1 0 158368 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_1466
timestamp 1698431365
transform 1 0 165536 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_1472
timestamp 1698431365
transform 1 0 166208 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_1536
timestamp 1698431365
transform 1 0 173376 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_1542
timestamp 1698431365
transform 1 0 174048 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_1606
timestamp 1698431365
transform 1 0 181216 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_1612
timestamp 1698431365
transform 1 0 181888 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_1676
timestamp 1698431365
transform 1 0 189056 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_1682
timestamp 1698431365
transform 1 0 189728 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_1746
timestamp 1698431365
transform 1 0 196896 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_1752
timestamp 1698431365
transform 1 0 197568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_1816
timestamp 1698431365
transform 1 0 204736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_1822
timestamp 1698431365
transform 1 0 205408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_1886
timestamp 1698431365
transform 1 0 212576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_1892
timestamp 1698431365
transform 1 0 213248 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_1924
timestamp 1698431365
transform 1 0 216832 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_1932
timestamp 1698431365
transform 1 0 217728 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_1936
timestamp 1698431365
transform 1 0 218176 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698431365
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698431365
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698431365
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698431365
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_317
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_381
timestamp 1698431365
transform 1 0 44016 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_387
timestamp 1698431365
transform 1 0 44688 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_451
timestamp 1698431365
transform 1 0 51856 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_457
timestamp 1698431365
transform 1 0 52528 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_521
timestamp 1698431365
transform 1 0 59696 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_527
timestamp 1698431365
transform 1 0 60368 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_591
timestamp 1698431365
transform 1 0 67536 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_597
timestamp 1698431365
transform 1 0 68208 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_661
timestamp 1698431365
transform 1 0 75376 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_667
timestamp 1698431365
transform 1 0 76048 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_731
timestamp 1698431365
transform 1 0 83216 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_737
timestamp 1698431365
transform 1 0 83888 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_801
timestamp 1698431365
transform 1 0 91056 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_807
timestamp 1698431365
transform 1 0 91728 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_871
timestamp 1698431365
transform 1 0 98896 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_877
timestamp 1698431365
transform 1 0 99568 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_941
timestamp 1698431365
transform 1 0 106736 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_947
timestamp 1698431365
transform 1 0 107408 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1011
timestamp 1698431365
transform 1 0 114576 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_1017
timestamp 1698431365
transform 1 0 115248 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1081
timestamp 1698431365
transform 1 0 122416 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_1087
timestamp 1698431365
transform 1 0 123088 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1151
timestamp 1698431365
transform 1 0 130256 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_1157
timestamp 1698431365
transform 1 0 130928 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1221
timestamp 1698431365
transform 1 0 138096 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_1227
timestamp 1698431365
transform 1 0 138768 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1231
timestamp 1698431365
transform 1 0 139216 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_1235
timestamp 1698431365
transform 1 0 139664 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_1238
timestamp 1698431365
transform 1 0 140000 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_1240
timestamp 1698431365
transform 1 0 140224 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_1253
timestamp 1698431365
transform 1 0 141680 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_1285
timestamp 1698431365
transform 1 0 145264 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_1293
timestamp 1698431365
transform 1 0 146160 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_1297
timestamp 1698431365
transform 1 0 146608 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1305
timestamp 1698431365
transform 1 0 147504 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_1309
timestamp 1698431365
transform 1 0 147952 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_1351
timestamp 1698431365
transform 1 0 152656 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1359
timestamp 1698431365
transform 1 0 153552 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_1367
timestamp 1698431365
transform 1 0 154448 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_1384
timestamp 1698431365
transform 1 0 156352 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_1386
timestamp 1698431365
transform 1 0 156576 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_1396
timestamp 1698431365
transform 1 0 157696 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_1400
timestamp 1698431365
transform 1 0 158144 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_1416
timestamp 1698431365
transform 1 0 159936 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_1424
timestamp 1698431365
transform 1 0 160832 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_1427
timestamp 1698431365
transform 1 0 161168 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_1437
timestamp 1698431365
transform 1 0 162288 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1501
timestamp 1698431365
transform 1 0 169456 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_1507
timestamp 1698431365
transform 1 0 170128 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1571
timestamp 1698431365
transform 1 0 177296 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_1577
timestamp 1698431365
transform 1 0 177968 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1641
timestamp 1698431365
transform 1 0 185136 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_1647
timestamp 1698431365
transform 1 0 185808 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1711
timestamp 1698431365
transform 1 0 192976 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_1717
timestamp 1698431365
transform 1 0 193648 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1781
timestamp 1698431365
transform 1 0 200816 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_1787
timestamp 1698431365
transform 1 0 201488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1851
timestamp 1698431365
transform 1 0 208656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_1857
timestamp 1698431365
transform 1 0 209328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_1921
timestamp 1698431365
transform 1 0 216496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_1927
timestamp 1698431365
transform 1 0 217168 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_1935
timestamp 1698431365
transform 1 0 218064 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_1937
timestamp 1698431365
transform 1 0 218288 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698431365
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698431365
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698431365
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698431365
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698431365
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_346
timestamp 1698431365
transform 1 0 40096 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_352
timestamp 1698431365
transform 1 0 40768 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_416
timestamp 1698431365
transform 1 0 47936 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_422
timestamp 1698431365
transform 1 0 48608 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_486
timestamp 1698431365
transform 1 0 55776 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_492
timestamp 1698431365
transform 1 0 56448 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_556
timestamp 1698431365
transform 1 0 63616 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_562
timestamp 1698431365
transform 1 0 64288 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_626
timestamp 1698431365
transform 1 0 71456 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_632
timestamp 1698431365
transform 1 0 72128 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_696
timestamp 1698431365
transform 1 0 79296 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_702
timestamp 1698431365
transform 1 0 79968 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_766
timestamp 1698431365
transform 1 0 87136 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_772
timestamp 1698431365
transform 1 0 87808 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_836
timestamp 1698431365
transform 1 0 94976 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_842
timestamp 1698431365
transform 1 0 95648 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_906
timestamp 1698431365
transform 1 0 102816 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_912
timestamp 1698431365
transform 1 0 103488 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_976
timestamp 1698431365
transform 1 0 110656 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_982
timestamp 1698431365
transform 1 0 111328 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_1046
timestamp 1698431365
transform 1 0 118496 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_1052
timestamp 1698431365
transform 1 0 119168 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_1116
timestamp 1698431365
transform 1 0 126336 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_1122
timestamp 1698431365
transform 1 0 127008 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_1186
timestamp 1698431365
transform 1 0 134176 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_1192
timestamp 1698431365
transform 1 0 134848 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_1256
timestamp 1698431365
transform 1 0 142016 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_1262
timestamp 1698431365
transform 1 0 142688 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_1294
timestamp 1698431365
transform 1 0 146272 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_1302
timestamp 1698431365
transform 1 0 147168 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_1306
timestamp 1698431365
transform 1 0 147616 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_1326
timestamp 1698431365
transform 1 0 149856 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_1332
timestamp 1698431365
transform 1 0 150528 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_1336
timestamp 1698431365
transform 1 0 150976 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_1345
timestamp 1698431365
transform 1 0 151984 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_1353
timestamp 1698431365
transform 1 0 152880 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_1362
timestamp 1698431365
transform 1 0 153888 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_1364
timestamp 1698431365
transform 1 0 154112 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_1397
timestamp 1698431365
transform 1 0 157808 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_1399
timestamp 1698431365
transform 1 0 158032 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_1402
timestamp 1698431365
transform 1 0 158368 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_1410
timestamp 1698431365
transform 1 0 159264 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_1414
timestamp 1698431365
transform 1 0 159712 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_1425
timestamp 1698431365
transform 1 0 160944 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_1441
timestamp 1698431365
transform 1 0 162736 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_1454
timestamp 1698431365
transform 1 0 164192 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_1458
timestamp 1698431365
transform 1 0 164640 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_1466
timestamp 1698431365
transform 1 0 165536 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_1472
timestamp 1698431365
transform 1 0 166208 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_1536
timestamp 1698431365
transform 1 0 173376 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_1542
timestamp 1698431365
transform 1 0 174048 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_1606
timestamp 1698431365
transform 1 0 181216 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_1612
timestamp 1698431365
transform 1 0 181888 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_1676
timestamp 1698431365
transform 1 0 189056 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_1682
timestamp 1698431365
transform 1 0 189728 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_1746
timestamp 1698431365
transform 1 0 196896 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_1752
timestamp 1698431365
transform 1 0 197568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_1816
timestamp 1698431365
transform 1 0 204736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_1822
timestamp 1698431365
transform 1 0 205408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_1886
timestamp 1698431365
transform 1 0 212576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_1892
timestamp 1698431365
transform 1 0 213248 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_1924
timestamp 1698431365
transform 1 0 216832 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_1932
timestamp 1698431365
transform 1 0 217728 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_1936
timestamp 1698431365
transform 1 0 218176 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698431365
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698431365
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698431365
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698431365
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698431365
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_317
timestamp 1698431365
transform 1 0 36848 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_381
timestamp 1698431365
transform 1 0 44016 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_387
timestamp 1698431365
transform 1 0 44688 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_451
timestamp 1698431365
transform 1 0 51856 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_457
timestamp 1698431365
transform 1 0 52528 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_521
timestamp 1698431365
transform 1 0 59696 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_527
timestamp 1698431365
transform 1 0 60368 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_591
timestamp 1698431365
transform 1 0 67536 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_597
timestamp 1698431365
transform 1 0 68208 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_661
timestamp 1698431365
transform 1 0 75376 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_667
timestamp 1698431365
transform 1 0 76048 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_731
timestamp 1698431365
transform 1 0 83216 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_737
timestamp 1698431365
transform 1 0 83888 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_801
timestamp 1698431365
transform 1 0 91056 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_807
timestamp 1698431365
transform 1 0 91728 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_871
timestamp 1698431365
transform 1 0 98896 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_877
timestamp 1698431365
transform 1 0 99568 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_941
timestamp 1698431365
transform 1 0 106736 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_947
timestamp 1698431365
transform 1 0 107408 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1011
timestamp 1698431365
transform 1 0 114576 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_1017
timestamp 1698431365
transform 1 0 115248 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1081
timestamp 1698431365
transform 1 0 122416 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_1087
timestamp 1698431365
transform 1 0 123088 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1151
timestamp 1698431365
transform 1 0 130256 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_1157
timestamp 1698431365
transform 1 0 130928 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1221
timestamp 1698431365
transform 1 0 138096 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_1227
timestamp 1698431365
transform 1 0 138768 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_1291
timestamp 1698431365
transform 1 0 145936 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_1297
timestamp 1698431365
transform 1 0 146608 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_1301
timestamp 1698431365
transform 1 0 147056 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_1318
timestamp 1698431365
transform 1 0 148960 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1322
timestamp 1698431365
transform 1 0 149408 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_1326
timestamp 1698431365
transform 1 0 149856 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_1333
timestamp 1698431365
transform 1 0 150640 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1367
timestamp 1698431365
transform 1 0 154448 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_1371
timestamp 1698431365
transform 1 0 154896 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1380
timestamp 1698431365
transform 1 0 155904 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_1393
timestamp 1698431365
transform 1 0 157360 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_1397
timestamp 1698431365
transform 1 0 157808 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1429
timestamp 1698431365
transform 1 0 161392 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_1433
timestamp 1698431365
transform 1 0 161840 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_1455
timestamp 1698431365
transform 1 0 164304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_1459
timestamp 1698431365
transform 1 0 164752 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_1491
timestamp 1698431365
transform 1 0 168336 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1499
timestamp 1698431365
transform 1 0 169232 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_1503
timestamp 1698431365
transform 1 0 169680 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_1507
timestamp 1698431365
transform 1 0 170128 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1571
timestamp 1698431365
transform 1 0 177296 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_1577
timestamp 1698431365
transform 1 0 177968 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1641
timestamp 1698431365
transform 1 0 185136 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_1647
timestamp 1698431365
transform 1 0 185808 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1711
timestamp 1698431365
transform 1 0 192976 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_1717
timestamp 1698431365
transform 1 0 193648 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1781
timestamp 1698431365
transform 1 0 200816 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_1787
timestamp 1698431365
transform 1 0 201488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1851
timestamp 1698431365
transform 1 0 208656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_1857
timestamp 1698431365
transform 1 0 209328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_1921
timestamp 1698431365
transform 1 0 216496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_1927
timestamp 1698431365
transform 1 0 217168 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_1935
timestamp 1698431365
transform 1 0 218064 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_1937
timestamp 1698431365
transform 1 0 218288 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698431365
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698431365
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698431365
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698431365
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698431365
transform 1 0 32928 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_346
timestamp 1698431365
transform 1 0 40096 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_352
timestamp 1698431365
transform 1 0 40768 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_416
timestamp 1698431365
transform 1 0 47936 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_422
timestamp 1698431365
transform 1 0 48608 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_486
timestamp 1698431365
transform 1 0 55776 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_492
timestamp 1698431365
transform 1 0 56448 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_556
timestamp 1698431365
transform 1 0 63616 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_562
timestamp 1698431365
transform 1 0 64288 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_626
timestamp 1698431365
transform 1 0 71456 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_632
timestamp 1698431365
transform 1 0 72128 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_696
timestamp 1698431365
transform 1 0 79296 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_702
timestamp 1698431365
transform 1 0 79968 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_766
timestamp 1698431365
transform 1 0 87136 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_772
timestamp 1698431365
transform 1 0 87808 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_836
timestamp 1698431365
transform 1 0 94976 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_842
timestamp 1698431365
transform 1 0 95648 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_906
timestamp 1698431365
transform 1 0 102816 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_912
timestamp 1698431365
transform 1 0 103488 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_976
timestamp 1698431365
transform 1 0 110656 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_982
timestamp 1698431365
transform 1 0 111328 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1046
timestamp 1698431365
transform 1 0 118496 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_1052
timestamp 1698431365
transform 1 0 119168 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1116
timestamp 1698431365
transform 1 0 126336 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_1122
timestamp 1698431365
transform 1 0 127008 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1186
timestamp 1698431365
transform 1 0 134176 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_1192
timestamp 1698431365
transform 1 0 134848 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1256
timestamp 1698431365
transform 1 0 142016 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_1262
timestamp 1698431365
transform 1 0 142688 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1326
timestamp 1698431365
transform 1 0 149856 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_1332
timestamp 1698431365
transform 1 0 150528 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_1364
timestamp 1698431365
transform 1 0 154112 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1372
timestamp 1698431365
transform 1 0 155008 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_1376
timestamp 1698431365
transform 1 0 155456 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_1378
timestamp 1698431365
transform 1 0 155680 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_1387
timestamp 1698431365
transform 1 0 156688 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1395
timestamp 1698431365
transform 1 0 157584 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_1399
timestamp 1698431365
transform 1 0 158032 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_1402
timestamp 1698431365
transform 1 0 158368 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_1434
timestamp 1698431365
transform 1 0 161952 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1442
timestamp 1698431365
transform 1 0 162848 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_1448
timestamp 1698431365
transform 1 0 163520 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1464
timestamp 1698431365
transform 1 0 165312 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_1468
timestamp 1698431365
transform 1 0 165760 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_1472
timestamp 1698431365
transform 1 0 166208 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1536
timestamp 1698431365
transform 1 0 173376 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_1542
timestamp 1698431365
transform 1 0 174048 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1606
timestamp 1698431365
transform 1 0 181216 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_1612
timestamp 1698431365
transform 1 0 181888 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1676
timestamp 1698431365
transform 1 0 189056 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_1682
timestamp 1698431365
transform 1 0 189728 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1746
timestamp 1698431365
transform 1 0 196896 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_1752
timestamp 1698431365
transform 1 0 197568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1816
timestamp 1698431365
transform 1 0 204736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_1822
timestamp 1698431365
transform 1 0 205408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1886
timestamp 1698431365
transform 1 0 212576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_1892
timestamp 1698431365
transform 1 0 213248 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_1924
timestamp 1698431365
transform 1 0 216832 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_1932
timestamp 1698431365
transform 1 0 217728 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_1936
timestamp 1698431365
transform 1 0 218176 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698431365
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698431365
transform 1 0 20496 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698431365
transform 1 0 28336 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698431365
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_317
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_381
timestamp 1698431365
transform 1 0 44016 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_387
timestamp 1698431365
transform 1 0 44688 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_451
timestamp 1698431365
transform 1 0 51856 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_457
timestamp 1698431365
transform 1 0 52528 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_521
timestamp 1698431365
transform 1 0 59696 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_527
timestamp 1698431365
transform 1 0 60368 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_591
timestamp 1698431365
transform 1 0 67536 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_597
timestamp 1698431365
transform 1 0 68208 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_661
timestamp 1698431365
transform 1 0 75376 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_667
timestamp 1698431365
transform 1 0 76048 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_731
timestamp 1698431365
transform 1 0 83216 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_737
timestamp 1698431365
transform 1 0 83888 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_801
timestamp 1698431365
transform 1 0 91056 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_807
timestamp 1698431365
transform 1 0 91728 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_871
timestamp 1698431365
transform 1 0 98896 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_877
timestamp 1698431365
transform 1 0 99568 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_941
timestamp 1698431365
transform 1 0 106736 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_947
timestamp 1698431365
transform 1 0 107408 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_1011
timestamp 1698431365
transform 1 0 114576 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_1017
timestamp 1698431365
transform 1 0 115248 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_1081
timestamp 1698431365
transform 1 0 122416 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_1087
timestamp 1698431365
transform 1 0 123088 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_1151
timestamp 1698431365
transform 1 0 130256 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_1157
timestamp 1698431365
transform 1 0 130928 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_1221
timestamp 1698431365
transform 1 0 138096 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_1227
timestamp 1698431365
transform 1 0 138768 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_1291
timestamp 1698431365
transform 1 0 145936 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_1297
timestamp 1698431365
transform 1 0 146608 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_1361
timestamp 1698431365
transform 1 0 153776 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_1367
timestamp 1698431365
transform 1 0 154448 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_1431
timestamp 1698431365
transform 1 0 161616 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_1437
timestamp 1698431365
transform 1 0 162288 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_1501
timestamp 1698431365
transform 1 0 169456 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_1507
timestamp 1698431365
transform 1 0 170128 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_1571
timestamp 1698431365
transform 1 0 177296 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_1577
timestamp 1698431365
transform 1 0 177968 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_1641
timestamp 1698431365
transform 1 0 185136 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_1647
timestamp 1698431365
transform 1 0 185808 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_1711
timestamp 1698431365
transform 1 0 192976 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_1717
timestamp 1698431365
transform 1 0 193648 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_1781
timestamp 1698431365
transform 1 0 200816 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_1787
timestamp 1698431365
transform 1 0 201488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_1851
timestamp 1698431365
transform 1 0 208656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_1857
timestamp 1698431365
transform 1 0 209328 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_1921
timestamp 1698431365
transform 1 0 216496 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_1927
timestamp 1698431365
transform 1 0 217168 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_1935
timestamp 1698431365
transform 1 0 218064 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_1937
timestamp 1698431365
transform 1 0 218288 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698431365
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698431365
transform 1 0 16576 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_206
timestamp 1698431365
transform 1 0 24416 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698431365
transform 1 0 32256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_346
timestamp 1698431365
transform 1 0 40096 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_352
timestamp 1698431365
transform 1 0 40768 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_416
timestamp 1698431365
transform 1 0 47936 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_422
timestamp 1698431365
transform 1 0 48608 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_486
timestamp 1698431365
transform 1 0 55776 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_492
timestamp 1698431365
transform 1 0 56448 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_556
timestamp 1698431365
transform 1 0 63616 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_562
timestamp 1698431365
transform 1 0 64288 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_626
timestamp 1698431365
transform 1 0 71456 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_632
timestamp 1698431365
transform 1 0 72128 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_696
timestamp 1698431365
transform 1 0 79296 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_702
timestamp 1698431365
transform 1 0 79968 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_766
timestamp 1698431365
transform 1 0 87136 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_772
timestamp 1698431365
transform 1 0 87808 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_836
timestamp 1698431365
transform 1 0 94976 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_842
timestamp 1698431365
transform 1 0 95648 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_906
timestamp 1698431365
transform 1 0 102816 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_912
timestamp 1698431365
transform 1 0 103488 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_976
timestamp 1698431365
transform 1 0 110656 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_982
timestamp 1698431365
transform 1 0 111328 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_1046
timestamp 1698431365
transform 1 0 118496 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_1052
timestamp 1698431365
transform 1 0 119168 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_1116
timestamp 1698431365
transform 1 0 126336 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_1122
timestamp 1698431365
transform 1 0 127008 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_1186
timestamp 1698431365
transform 1 0 134176 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_1192
timestamp 1698431365
transform 1 0 134848 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_1256
timestamp 1698431365
transform 1 0 142016 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_1262
timestamp 1698431365
transform 1 0 142688 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_1326
timestamp 1698431365
transform 1 0 149856 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_1332
timestamp 1698431365
transform 1 0 150528 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_1396
timestamp 1698431365
transform 1 0 157696 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_1402
timestamp 1698431365
transform 1 0 158368 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_1466
timestamp 1698431365
transform 1 0 165536 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_1472
timestamp 1698431365
transform 1 0 166208 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_1536
timestamp 1698431365
transform 1 0 173376 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_1542
timestamp 1698431365
transform 1 0 174048 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_1606
timestamp 1698431365
transform 1 0 181216 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_1612
timestamp 1698431365
transform 1 0 181888 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_1676
timestamp 1698431365
transform 1 0 189056 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_1682
timestamp 1698431365
transform 1 0 189728 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_1746
timestamp 1698431365
transform 1 0 196896 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_1752
timestamp 1698431365
transform 1 0 197568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_1816
timestamp 1698431365
transform 1 0 204736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_1822
timestamp 1698431365
transform 1 0 205408 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_1886
timestamp 1698431365
transform 1 0 212576 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_1892
timestamp 1698431365
transform 1 0 213248 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_1924
timestamp 1698431365
transform 1 0 216832 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_1932
timestamp 1698431365
transform 1 0 217728 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_1936
timestamp 1698431365
transform 1 0 218176 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698431365
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_171
timestamp 1698431365
transform 1 0 20496 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_177
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_241
timestamp 1698431365
transform 1 0 28336 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698431365
transform 1 0 36176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_317
timestamp 1698431365
transform 1 0 36848 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_381
timestamp 1698431365
transform 1 0 44016 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_387
timestamp 1698431365
transform 1 0 44688 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_451
timestamp 1698431365
transform 1 0 51856 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_457
timestamp 1698431365
transform 1 0 52528 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_521
timestamp 1698431365
transform 1 0 59696 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_527
timestamp 1698431365
transform 1 0 60368 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_591
timestamp 1698431365
transform 1 0 67536 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_597
timestamp 1698431365
transform 1 0 68208 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_661
timestamp 1698431365
transform 1 0 75376 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_667
timestamp 1698431365
transform 1 0 76048 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_731
timestamp 1698431365
transform 1 0 83216 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_737
timestamp 1698431365
transform 1 0 83888 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_801
timestamp 1698431365
transform 1 0 91056 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_807
timestamp 1698431365
transform 1 0 91728 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_871
timestamp 1698431365
transform 1 0 98896 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_877
timestamp 1698431365
transform 1 0 99568 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_941
timestamp 1698431365
transform 1 0 106736 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_947
timestamp 1698431365
transform 1 0 107408 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1011
timestamp 1698431365
transform 1 0 114576 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_1017
timestamp 1698431365
transform 1 0 115248 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1081
timestamp 1698431365
transform 1 0 122416 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_1087
timestamp 1698431365
transform 1 0 123088 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1151
timestamp 1698431365
transform 1 0 130256 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_1157
timestamp 1698431365
transform 1 0 130928 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1221
timestamp 1698431365
transform 1 0 138096 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_1227
timestamp 1698431365
transform 1 0 138768 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1291
timestamp 1698431365
transform 1 0 145936 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_1297
timestamp 1698431365
transform 1 0 146608 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1361
timestamp 1698431365
transform 1 0 153776 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_1367
timestamp 1698431365
transform 1 0 154448 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1431
timestamp 1698431365
transform 1 0 161616 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_1437
timestamp 1698431365
transform 1 0 162288 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1501
timestamp 1698431365
transform 1 0 169456 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_1507
timestamp 1698431365
transform 1 0 170128 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1571
timestamp 1698431365
transform 1 0 177296 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_1577
timestamp 1698431365
transform 1 0 177968 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1641
timestamp 1698431365
transform 1 0 185136 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_1647
timestamp 1698431365
transform 1 0 185808 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1711
timestamp 1698431365
transform 1 0 192976 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_1717
timestamp 1698431365
transform 1 0 193648 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1781
timestamp 1698431365
transform 1 0 200816 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_1787
timestamp 1698431365
transform 1 0 201488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1851
timestamp 1698431365
transform 1 0 208656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_1857
timestamp 1698431365
transform 1 0 209328 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_1921
timestamp 1698431365
transform 1 0 216496 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_1927
timestamp 1698431365
transform 1 0 217168 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_1935
timestamp 1698431365
transform 1 0 218064 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_1937
timestamp 1698431365
transform 1 0 218288 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698431365
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_72
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_136
timestamp 1698431365
transform 1 0 16576 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_142
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_206
timestamp 1698431365
transform 1 0 24416 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_212
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_276
timestamp 1698431365
transform 1 0 32256 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698431365
transform 1 0 32928 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_346
timestamp 1698431365
transform 1 0 40096 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_352
timestamp 1698431365
transform 1 0 40768 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_416
timestamp 1698431365
transform 1 0 47936 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_422
timestamp 1698431365
transform 1 0 48608 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_486
timestamp 1698431365
transform 1 0 55776 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_492
timestamp 1698431365
transform 1 0 56448 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_556
timestamp 1698431365
transform 1 0 63616 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_562
timestamp 1698431365
transform 1 0 64288 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_626
timestamp 1698431365
transform 1 0 71456 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_632
timestamp 1698431365
transform 1 0 72128 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_696
timestamp 1698431365
transform 1 0 79296 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_702
timestamp 1698431365
transform 1 0 79968 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_766
timestamp 1698431365
transform 1 0 87136 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_772
timestamp 1698431365
transform 1 0 87808 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_836
timestamp 1698431365
transform 1 0 94976 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_842
timestamp 1698431365
transform 1 0 95648 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_906
timestamp 1698431365
transform 1 0 102816 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_912
timestamp 1698431365
transform 1 0 103488 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_976
timestamp 1698431365
transform 1 0 110656 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_982
timestamp 1698431365
transform 1 0 111328 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_1046
timestamp 1698431365
transform 1 0 118496 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_1052
timestamp 1698431365
transform 1 0 119168 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_1116
timestamp 1698431365
transform 1 0 126336 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_1122
timestamp 1698431365
transform 1 0 127008 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_1186
timestamp 1698431365
transform 1 0 134176 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_1192
timestamp 1698431365
transform 1 0 134848 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_1256
timestamp 1698431365
transform 1 0 142016 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_1262
timestamp 1698431365
transform 1 0 142688 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_1326
timestamp 1698431365
transform 1 0 149856 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_1332
timestamp 1698431365
transform 1 0 150528 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_1396
timestamp 1698431365
transform 1 0 157696 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_1402
timestamp 1698431365
transform 1 0 158368 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_1466
timestamp 1698431365
transform 1 0 165536 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_1472
timestamp 1698431365
transform 1 0 166208 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_1536
timestamp 1698431365
transform 1 0 173376 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_1542
timestamp 1698431365
transform 1 0 174048 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_1606
timestamp 1698431365
transform 1 0 181216 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_1612
timestamp 1698431365
transform 1 0 181888 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_1676
timestamp 1698431365
transform 1 0 189056 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_1682
timestamp 1698431365
transform 1 0 189728 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_1746
timestamp 1698431365
transform 1 0 196896 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_1752
timestamp 1698431365
transform 1 0 197568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_1816
timestamp 1698431365
transform 1 0 204736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_1822
timestamp 1698431365
transform 1 0 205408 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_1886
timestamp 1698431365
transform 1 0 212576 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_1892
timestamp 1698431365
transform 1 0 213248 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_1924
timestamp 1698431365
transform 1 0 216832 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_1932
timestamp 1698431365
transform 1 0 217728 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_1936
timestamp 1698431365
transform 1 0 218176 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698431365
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698431365
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_107
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_171
timestamp 1698431365
transform 1 0 20496 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_177
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_241
timestamp 1698431365
transform 1 0 28336 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698431365
transform 1 0 36176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_317
timestamp 1698431365
transform 1 0 36848 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_381
timestamp 1698431365
transform 1 0 44016 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_387
timestamp 1698431365
transform 1 0 44688 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_451
timestamp 1698431365
transform 1 0 51856 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_457
timestamp 1698431365
transform 1 0 52528 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_521
timestamp 1698431365
transform 1 0 59696 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_527
timestamp 1698431365
transform 1 0 60368 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_591
timestamp 1698431365
transform 1 0 67536 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_597
timestamp 1698431365
transform 1 0 68208 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_661
timestamp 1698431365
transform 1 0 75376 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_667
timestamp 1698431365
transform 1 0 76048 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_731
timestamp 1698431365
transform 1 0 83216 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_737
timestamp 1698431365
transform 1 0 83888 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_801
timestamp 1698431365
transform 1 0 91056 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_807
timestamp 1698431365
transform 1 0 91728 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_871
timestamp 1698431365
transform 1 0 98896 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_877
timestamp 1698431365
transform 1 0 99568 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_941
timestamp 1698431365
transform 1 0 106736 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_947
timestamp 1698431365
transform 1 0 107408 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1011
timestamp 1698431365
transform 1 0 114576 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_1017
timestamp 1698431365
transform 1 0 115248 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1081
timestamp 1698431365
transform 1 0 122416 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_1087
timestamp 1698431365
transform 1 0 123088 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1151
timestamp 1698431365
transform 1 0 130256 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_1157
timestamp 1698431365
transform 1 0 130928 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1221
timestamp 1698431365
transform 1 0 138096 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_1227
timestamp 1698431365
transform 1 0 138768 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1291
timestamp 1698431365
transform 1 0 145936 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_1297
timestamp 1698431365
transform 1 0 146608 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1361
timestamp 1698431365
transform 1 0 153776 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_1367
timestamp 1698431365
transform 1 0 154448 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1431
timestamp 1698431365
transform 1 0 161616 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_1437
timestamp 1698431365
transform 1 0 162288 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1501
timestamp 1698431365
transform 1 0 169456 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_1507
timestamp 1698431365
transform 1 0 170128 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1571
timestamp 1698431365
transform 1 0 177296 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_1577
timestamp 1698431365
transform 1 0 177968 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1641
timestamp 1698431365
transform 1 0 185136 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_1647
timestamp 1698431365
transform 1 0 185808 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1711
timestamp 1698431365
transform 1 0 192976 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_1717
timestamp 1698431365
transform 1 0 193648 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1781
timestamp 1698431365
transform 1 0 200816 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_1787
timestamp 1698431365
transform 1 0 201488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1851
timestamp 1698431365
transform 1 0 208656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_1857
timestamp 1698431365
transform 1 0 209328 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_1921
timestamp 1698431365
transform 1 0 216496 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_1927
timestamp 1698431365
transform 1 0 217168 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_1935
timestamp 1698431365
transform 1 0 218064 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_1937
timestamp 1698431365
transform 1 0 218288 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698431365
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_72
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_136
timestamp 1698431365
transform 1 0 16576 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_142
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_206
timestamp 1698431365
transform 1 0 24416 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_212
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_276
timestamp 1698431365
transform 1 0 32256 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_282
timestamp 1698431365
transform 1 0 32928 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_346
timestamp 1698431365
transform 1 0 40096 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_352
timestamp 1698431365
transform 1 0 40768 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_416
timestamp 1698431365
transform 1 0 47936 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_422
timestamp 1698431365
transform 1 0 48608 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_486
timestamp 1698431365
transform 1 0 55776 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_492
timestamp 1698431365
transform 1 0 56448 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_556
timestamp 1698431365
transform 1 0 63616 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_562
timestamp 1698431365
transform 1 0 64288 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_626
timestamp 1698431365
transform 1 0 71456 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_632
timestamp 1698431365
transform 1 0 72128 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_696
timestamp 1698431365
transform 1 0 79296 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_702
timestamp 1698431365
transform 1 0 79968 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_766
timestamp 1698431365
transform 1 0 87136 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_772
timestamp 1698431365
transform 1 0 87808 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_836
timestamp 1698431365
transform 1 0 94976 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_842
timestamp 1698431365
transform 1 0 95648 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_906
timestamp 1698431365
transform 1 0 102816 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_912
timestamp 1698431365
transform 1 0 103488 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_976
timestamp 1698431365
transform 1 0 110656 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_982
timestamp 1698431365
transform 1 0 111328 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_1046
timestamp 1698431365
transform 1 0 118496 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_1052
timestamp 1698431365
transform 1 0 119168 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_1116
timestamp 1698431365
transform 1 0 126336 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_1122
timestamp 1698431365
transform 1 0 127008 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_1186
timestamp 1698431365
transform 1 0 134176 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_1192
timestamp 1698431365
transform 1 0 134848 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_1256
timestamp 1698431365
transform 1 0 142016 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_1262
timestamp 1698431365
transform 1 0 142688 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_1326
timestamp 1698431365
transform 1 0 149856 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_1332
timestamp 1698431365
transform 1 0 150528 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_1396
timestamp 1698431365
transform 1 0 157696 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_1402
timestamp 1698431365
transform 1 0 158368 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_1466
timestamp 1698431365
transform 1 0 165536 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_1472
timestamp 1698431365
transform 1 0 166208 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_1536
timestamp 1698431365
transform 1 0 173376 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_1542
timestamp 1698431365
transform 1 0 174048 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_1606
timestamp 1698431365
transform 1 0 181216 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_1612
timestamp 1698431365
transform 1 0 181888 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_1676
timestamp 1698431365
transform 1 0 189056 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_1682
timestamp 1698431365
transform 1 0 189728 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_1746
timestamp 1698431365
transform 1 0 196896 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_1752
timestamp 1698431365
transform 1 0 197568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_1816
timestamp 1698431365
transform 1 0 204736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_1822
timestamp 1698431365
transform 1 0 205408 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_1886
timestamp 1698431365
transform 1 0 212576 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_1892
timestamp 1698431365
transform 1 0 213248 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_1924
timestamp 1698431365
transform 1 0 216832 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_1932
timestamp 1698431365
transform 1 0 217728 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_1936
timestamp 1698431365
transform 1 0 218176 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698431365
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698431365
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_107
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_171
timestamp 1698431365
transform 1 0 20496 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_177
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_241
timestamp 1698431365
transform 1 0 28336 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698431365
transform 1 0 36176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_317
timestamp 1698431365
transform 1 0 36848 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_381
timestamp 1698431365
transform 1 0 44016 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_387
timestamp 1698431365
transform 1 0 44688 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_451
timestamp 1698431365
transform 1 0 51856 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_457
timestamp 1698431365
transform 1 0 52528 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_521
timestamp 1698431365
transform 1 0 59696 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_527
timestamp 1698431365
transform 1 0 60368 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_591
timestamp 1698431365
transform 1 0 67536 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_597
timestamp 1698431365
transform 1 0 68208 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_661
timestamp 1698431365
transform 1 0 75376 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_667
timestamp 1698431365
transform 1 0 76048 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_731
timestamp 1698431365
transform 1 0 83216 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_737
timestamp 1698431365
transform 1 0 83888 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_801
timestamp 1698431365
transform 1 0 91056 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_807
timestamp 1698431365
transform 1 0 91728 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_871
timestamp 1698431365
transform 1 0 98896 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_877
timestamp 1698431365
transform 1 0 99568 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_941
timestamp 1698431365
transform 1 0 106736 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_947
timestamp 1698431365
transform 1 0 107408 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_1011
timestamp 1698431365
transform 1 0 114576 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_1017
timestamp 1698431365
transform 1 0 115248 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_1081
timestamp 1698431365
transform 1 0 122416 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_1087
timestamp 1698431365
transform 1 0 123088 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_1151
timestamp 1698431365
transform 1 0 130256 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_1157
timestamp 1698431365
transform 1 0 130928 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_1221
timestamp 1698431365
transform 1 0 138096 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_1227
timestamp 1698431365
transform 1 0 138768 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_1291
timestamp 1698431365
transform 1 0 145936 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_1297
timestamp 1698431365
transform 1 0 146608 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_1361
timestamp 1698431365
transform 1 0 153776 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_1367
timestamp 1698431365
transform 1 0 154448 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_1431
timestamp 1698431365
transform 1 0 161616 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_1437
timestamp 1698431365
transform 1 0 162288 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_1501
timestamp 1698431365
transform 1 0 169456 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_1507
timestamp 1698431365
transform 1 0 170128 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_1571
timestamp 1698431365
transform 1 0 177296 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_1577
timestamp 1698431365
transform 1 0 177968 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_1641
timestamp 1698431365
transform 1 0 185136 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_1647
timestamp 1698431365
transform 1 0 185808 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_1711
timestamp 1698431365
transform 1 0 192976 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_1717
timestamp 1698431365
transform 1 0 193648 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_1781
timestamp 1698431365
transform 1 0 200816 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_1787
timestamp 1698431365
transform 1 0 201488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_1851
timestamp 1698431365
transform 1 0 208656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_1857
timestamp 1698431365
transform 1 0 209328 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_1921
timestamp 1698431365
transform 1 0 216496 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_1927
timestamp 1698431365
transform 1 0 217168 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_1935
timestamp 1698431365
transform 1 0 218064 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_1937
timestamp 1698431365
transform 1 0 218288 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698431365
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_136
timestamp 1698431365
transform 1 0 16576 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_206
timestamp 1698431365
transform 1 0 24416 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_212
timestamp 1698431365
transform 1 0 25088 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_276
timestamp 1698431365
transform 1 0 32256 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_282
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_346
timestamp 1698431365
transform 1 0 40096 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_352
timestamp 1698431365
transform 1 0 40768 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_416
timestamp 1698431365
transform 1 0 47936 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_422
timestamp 1698431365
transform 1 0 48608 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_486
timestamp 1698431365
transform 1 0 55776 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_492
timestamp 1698431365
transform 1 0 56448 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_556
timestamp 1698431365
transform 1 0 63616 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_562
timestamp 1698431365
transform 1 0 64288 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_626
timestamp 1698431365
transform 1 0 71456 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_632
timestamp 1698431365
transform 1 0 72128 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_696
timestamp 1698431365
transform 1 0 79296 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_702
timestamp 1698431365
transform 1 0 79968 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_766
timestamp 1698431365
transform 1 0 87136 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_772
timestamp 1698431365
transform 1 0 87808 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_836
timestamp 1698431365
transform 1 0 94976 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_842
timestamp 1698431365
transform 1 0 95648 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_906
timestamp 1698431365
transform 1 0 102816 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_912
timestamp 1698431365
transform 1 0 103488 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_976
timestamp 1698431365
transform 1 0 110656 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_982
timestamp 1698431365
transform 1 0 111328 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_1046
timestamp 1698431365
transform 1 0 118496 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_1052
timestamp 1698431365
transform 1 0 119168 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_1116
timestamp 1698431365
transform 1 0 126336 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_1122
timestamp 1698431365
transform 1 0 127008 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_1186
timestamp 1698431365
transform 1 0 134176 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_1192
timestamp 1698431365
transform 1 0 134848 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_1256
timestamp 1698431365
transform 1 0 142016 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_1262
timestamp 1698431365
transform 1 0 142688 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_1326
timestamp 1698431365
transform 1 0 149856 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_1332
timestamp 1698431365
transform 1 0 150528 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_1396
timestamp 1698431365
transform 1 0 157696 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_1402
timestamp 1698431365
transform 1 0 158368 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_1466
timestamp 1698431365
transform 1 0 165536 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_1472
timestamp 1698431365
transform 1 0 166208 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_1536
timestamp 1698431365
transform 1 0 173376 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_1542
timestamp 1698431365
transform 1 0 174048 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_1606
timestamp 1698431365
transform 1 0 181216 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_1612
timestamp 1698431365
transform 1 0 181888 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_1676
timestamp 1698431365
transform 1 0 189056 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_1682
timestamp 1698431365
transform 1 0 189728 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_1746
timestamp 1698431365
transform 1 0 196896 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_1752
timestamp 1698431365
transform 1 0 197568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_1816
timestamp 1698431365
transform 1 0 204736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_1822
timestamp 1698431365
transform 1 0 205408 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_1886
timestamp 1698431365
transform 1 0 212576 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_1892
timestamp 1698431365
transform 1 0 213248 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_1924
timestamp 1698431365
transform 1 0 216832 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_1932
timestamp 1698431365
transform 1 0 217728 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_1936
timestamp 1698431365
transform 1 0 218176 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698431365
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698431365
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_107
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_171
timestamp 1698431365
transform 1 0 20496 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_177
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_241
timestamp 1698431365
transform 1 0 28336 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698431365
transform 1 0 36176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_317
timestamp 1698431365
transform 1 0 36848 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_381
timestamp 1698431365
transform 1 0 44016 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_387
timestamp 1698431365
transform 1 0 44688 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_451
timestamp 1698431365
transform 1 0 51856 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_457
timestamp 1698431365
transform 1 0 52528 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_521
timestamp 1698431365
transform 1 0 59696 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_527
timestamp 1698431365
transform 1 0 60368 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_591
timestamp 1698431365
transform 1 0 67536 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_597
timestamp 1698431365
transform 1 0 68208 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_661
timestamp 1698431365
transform 1 0 75376 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_667
timestamp 1698431365
transform 1 0 76048 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_731
timestamp 1698431365
transform 1 0 83216 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_737
timestamp 1698431365
transform 1 0 83888 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_801
timestamp 1698431365
transform 1 0 91056 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_807
timestamp 1698431365
transform 1 0 91728 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_871
timestamp 1698431365
transform 1 0 98896 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_877
timestamp 1698431365
transform 1 0 99568 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_941
timestamp 1698431365
transform 1 0 106736 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_947
timestamp 1698431365
transform 1 0 107408 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_1011
timestamp 1698431365
transform 1 0 114576 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_1017
timestamp 1698431365
transform 1 0 115248 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_1081
timestamp 1698431365
transform 1 0 122416 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_1087
timestamp 1698431365
transform 1 0 123088 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_1151
timestamp 1698431365
transform 1 0 130256 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_1157
timestamp 1698431365
transform 1 0 130928 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_1221
timestamp 1698431365
transform 1 0 138096 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_1227
timestamp 1698431365
transform 1 0 138768 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_1291
timestamp 1698431365
transform 1 0 145936 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_1297
timestamp 1698431365
transform 1 0 146608 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_1361
timestamp 1698431365
transform 1 0 153776 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_1367
timestamp 1698431365
transform 1 0 154448 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_1431
timestamp 1698431365
transform 1 0 161616 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_1437
timestamp 1698431365
transform 1 0 162288 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_1501
timestamp 1698431365
transform 1 0 169456 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_1507
timestamp 1698431365
transform 1 0 170128 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_1571
timestamp 1698431365
transform 1 0 177296 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_1577
timestamp 1698431365
transform 1 0 177968 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_1641
timestamp 1698431365
transform 1 0 185136 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_1647
timestamp 1698431365
transform 1 0 185808 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_1711
timestamp 1698431365
transform 1 0 192976 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_1717
timestamp 1698431365
transform 1 0 193648 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_1781
timestamp 1698431365
transform 1 0 200816 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_1787
timestamp 1698431365
transform 1 0 201488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_1851
timestamp 1698431365
transform 1 0 208656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_1857
timestamp 1698431365
transform 1 0 209328 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_1921
timestamp 1698431365
transform 1 0 216496 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_1927
timestamp 1698431365
transform 1 0 217168 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_1935
timestamp 1698431365
transform 1 0 218064 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_1937
timestamp 1698431365
transform 1 0 218288 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698431365
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_72
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_136
timestamp 1698431365
transform 1 0 16576 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_142
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_206
timestamp 1698431365
transform 1 0 24416 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_212
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_276
timestamp 1698431365
transform 1 0 32256 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_282
timestamp 1698431365
transform 1 0 32928 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_346
timestamp 1698431365
transform 1 0 40096 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_352
timestamp 1698431365
transform 1 0 40768 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_416
timestamp 1698431365
transform 1 0 47936 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_422
timestamp 1698431365
transform 1 0 48608 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_486
timestamp 1698431365
transform 1 0 55776 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_492
timestamp 1698431365
transform 1 0 56448 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_556
timestamp 1698431365
transform 1 0 63616 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_562
timestamp 1698431365
transform 1 0 64288 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_626
timestamp 1698431365
transform 1 0 71456 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_632
timestamp 1698431365
transform 1 0 72128 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_696
timestamp 1698431365
transform 1 0 79296 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_702
timestamp 1698431365
transform 1 0 79968 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_766
timestamp 1698431365
transform 1 0 87136 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_772
timestamp 1698431365
transform 1 0 87808 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_836
timestamp 1698431365
transform 1 0 94976 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_842
timestamp 1698431365
transform 1 0 95648 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_906
timestamp 1698431365
transform 1 0 102816 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_912
timestamp 1698431365
transform 1 0 103488 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_976
timestamp 1698431365
transform 1 0 110656 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_982
timestamp 1698431365
transform 1 0 111328 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_1046
timestamp 1698431365
transform 1 0 118496 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_1052
timestamp 1698431365
transform 1 0 119168 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_1116
timestamp 1698431365
transform 1 0 126336 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_1122
timestamp 1698431365
transform 1 0 127008 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_1186
timestamp 1698431365
transform 1 0 134176 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_1192
timestamp 1698431365
transform 1 0 134848 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_1256
timestamp 1698431365
transform 1 0 142016 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_1262
timestamp 1698431365
transform 1 0 142688 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_1326
timestamp 1698431365
transform 1 0 149856 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_1332
timestamp 1698431365
transform 1 0 150528 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_1396
timestamp 1698431365
transform 1 0 157696 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_1402
timestamp 1698431365
transform 1 0 158368 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_1466
timestamp 1698431365
transform 1 0 165536 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_1472
timestamp 1698431365
transform 1 0 166208 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_1536
timestamp 1698431365
transform 1 0 173376 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_1542
timestamp 1698431365
transform 1 0 174048 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_1606
timestamp 1698431365
transform 1 0 181216 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_1612
timestamp 1698431365
transform 1 0 181888 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_1676
timestamp 1698431365
transform 1 0 189056 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_1682
timestamp 1698431365
transform 1 0 189728 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_1746
timestamp 1698431365
transform 1 0 196896 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_1752
timestamp 1698431365
transform 1 0 197568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_1816
timestamp 1698431365
transform 1 0 204736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_1822
timestamp 1698431365
transform 1 0 205408 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_1886
timestamp 1698431365
transform 1 0 212576 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_1892
timestamp 1698431365
transform 1 0 213248 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_1924
timestamp 1698431365
transform 1 0 216832 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_1932
timestamp 1698431365
transform 1 0 217728 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_1936
timestamp 1698431365
transform 1 0 218176 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698431365
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698431365
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_107
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_171
timestamp 1698431365
transform 1 0 20496 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_177
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_241
timestamp 1698431365
transform 1 0 28336 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698431365
transform 1 0 29008 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698431365
transform 1 0 36176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_317
timestamp 1698431365
transform 1 0 36848 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_381
timestamp 1698431365
transform 1 0 44016 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_387
timestamp 1698431365
transform 1 0 44688 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_451
timestamp 1698431365
transform 1 0 51856 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_457
timestamp 1698431365
transform 1 0 52528 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_521
timestamp 1698431365
transform 1 0 59696 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_527
timestamp 1698431365
transform 1 0 60368 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_591
timestamp 1698431365
transform 1 0 67536 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_597
timestamp 1698431365
transform 1 0 68208 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_661
timestamp 1698431365
transform 1 0 75376 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_667
timestamp 1698431365
transform 1 0 76048 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_731
timestamp 1698431365
transform 1 0 83216 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_737
timestamp 1698431365
transform 1 0 83888 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_801
timestamp 1698431365
transform 1 0 91056 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_807
timestamp 1698431365
transform 1 0 91728 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_871
timestamp 1698431365
transform 1 0 98896 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_877
timestamp 1698431365
transform 1 0 99568 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_941
timestamp 1698431365
transform 1 0 106736 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_947
timestamp 1698431365
transform 1 0 107408 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_1011
timestamp 1698431365
transform 1 0 114576 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_1017
timestamp 1698431365
transform 1 0 115248 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_1081
timestamp 1698431365
transform 1 0 122416 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_1087
timestamp 1698431365
transform 1 0 123088 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_1151
timestamp 1698431365
transform 1 0 130256 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_1157
timestamp 1698431365
transform 1 0 130928 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_1221
timestamp 1698431365
transform 1 0 138096 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_1227
timestamp 1698431365
transform 1 0 138768 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_1291
timestamp 1698431365
transform 1 0 145936 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_1297
timestamp 1698431365
transform 1 0 146608 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_1361
timestamp 1698431365
transform 1 0 153776 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_1367
timestamp 1698431365
transform 1 0 154448 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_1431
timestamp 1698431365
transform 1 0 161616 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_1437
timestamp 1698431365
transform 1 0 162288 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_1501
timestamp 1698431365
transform 1 0 169456 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_1507
timestamp 1698431365
transform 1 0 170128 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_1571
timestamp 1698431365
transform 1 0 177296 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_1577
timestamp 1698431365
transform 1 0 177968 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_1641
timestamp 1698431365
transform 1 0 185136 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_1647
timestamp 1698431365
transform 1 0 185808 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_1711
timestamp 1698431365
transform 1 0 192976 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_1717
timestamp 1698431365
transform 1 0 193648 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_1781
timestamp 1698431365
transform 1 0 200816 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_1787
timestamp 1698431365
transform 1 0 201488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_1851
timestamp 1698431365
transform 1 0 208656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_1857
timestamp 1698431365
transform 1 0 209328 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_1921
timestamp 1698431365
transform 1 0 216496 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_1927
timestamp 1698431365
transform 1 0 217168 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_1935
timestamp 1698431365
transform 1 0 218064 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_1937
timestamp 1698431365
transform 1 0 218288 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698431365
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_136
timestamp 1698431365
transform 1 0 16576 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_142
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_206
timestamp 1698431365
transform 1 0 24416 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_212
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_276
timestamp 1698431365
transform 1 0 32256 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_282
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_346
timestamp 1698431365
transform 1 0 40096 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_352
timestamp 1698431365
transform 1 0 40768 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_416
timestamp 1698431365
transform 1 0 47936 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_422
timestamp 1698431365
transform 1 0 48608 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_486
timestamp 1698431365
transform 1 0 55776 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_492
timestamp 1698431365
transform 1 0 56448 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_556
timestamp 1698431365
transform 1 0 63616 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_562
timestamp 1698431365
transform 1 0 64288 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_626
timestamp 1698431365
transform 1 0 71456 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_632
timestamp 1698431365
transform 1 0 72128 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_696
timestamp 1698431365
transform 1 0 79296 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_702
timestamp 1698431365
transform 1 0 79968 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_766
timestamp 1698431365
transform 1 0 87136 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_772
timestamp 1698431365
transform 1 0 87808 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_836
timestamp 1698431365
transform 1 0 94976 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_842
timestamp 1698431365
transform 1 0 95648 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_906
timestamp 1698431365
transform 1 0 102816 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_912
timestamp 1698431365
transform 1 0 103488 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_976
timestamp 1698431365
transform 1 0 110656 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_982
timestamp 1698431365
transform 1 0 111328 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_1046
timestamp 1698431365
transform 1 0 118496 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_1052
timestamp 1698431365
transform 1 0 119168 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_1116
timestamp 1698431365
transform 1 0 126336 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_1122
timestamp 1698431365
transform 1 0 127008 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_1186
timestamp 1698431365
transform 1 0 134176 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_1192
timestamp 1698431365
transform 1 0 134848 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_1256
timestamp 1698431365
transform 1 0 142016 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_1262
timestamp 1698431365
transform 1 0 142688 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_1326
timestamp 1698431365
transform 1 0 149856 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_1332
timestamp 1698431365
transform 1 0 150528 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_1396
timestamp 1698431365
transform 1 0 157696 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_1402
timestamp 1698431365
transform 1 0 158368 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_1466
timestamp 1698431365
transform 1 0 165536 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_1472
timestamp 1698431365
transform 1 0 166208 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_1536
timestamp 1698431365
transform 1 0 173376 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_1542
timestamp 1698431365
transform 1 0 174048 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_1606
timestamp 1698431365
transform 1 0 181216 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_1612
timestamp 1698431365
transform 1 0 181888 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_1676
timestamp 1698431365
transform 1 0 189056 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_1682
timestamp 1698431365
transform 1 0 189728 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_1746
timestamp 1698431365
transform 1 0 196896 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_1752
timestamp 1698431365
transform 1 0 197568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_1816
timestamp 1698431365
transform 1 0 204736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_1822
timestamp 1698431365
transform 1 0 205408 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_1886
timestamp 1698431365
transform 1 0 212576 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_1892
timestamp 1698431365
transform 1 0 213248 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_1924
timestamp 1698431365
transform 1 0 216832 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_1932
timestamp 1698431365
transform 1 0 217728 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_1936
timestamp 1698431365
transform 1 0 218176 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698431365
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698431365
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_107
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_171
timestamp 1698431365
transform 1 0 20496 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_177
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_241
timestamp 1698431365
transform 1 0 28336 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698431365
transform 1 0 29008 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698431365
transform 1 0 36176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_317
timestamp 1698431365
transform 1 0 36848 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_381
timestamp 1698431365
transform 1 0 44016 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_387
timestamp 1698431365
transform 1 0 44688 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_451
timestamp 1698431365
transform 1 0 51856 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_457
timestamp 1698431365
transform 1 0 52528 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_521
timestamp 1698431365
transform 1 0 59696 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_527
timestamp 1698431365
transform 1 0 60368 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_591
timestamp 1698431365
transform 1 0 67536 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_597
timestamp 1698431365
transform 1 0 68208 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_661
timestamp 1698431365
transform 1 0 75376 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_667
timestamp 1698431365
transform 1 0 76048 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_731
timestamp 1698431365
transform 1 0 83216 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_737
timestamp 1698431365
transform 1 0 83888 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_801
timestamp 1698431365
transform 1 0 91056 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_807
timestamp 1698431365
transform 1 0 91728 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_871
timestamp 1698431365
transform 1 0 98896 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_877
timestamp 1698431365
transform 1 0 99568 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_941
timestamp 1698431365
transform 1 0 106736 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_947
timestamp 1698431365
transform 1 0 107408 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_1011
timestamp 1698431365
transform 1 0 114576 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_1017
timestamp 1698431365
transform 1 0 115248 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_1081
timestamp 1698431365
transform 1 0 122416 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_1087
timestamp 1698431365
transform 1 0 123088 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_1151
timestamp 1698431365
transform 1 0 130256 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_1157
timestamp 1698431365
transform 1 0 130928 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_1221
timestamp 1698431365
transform 1 0 138096 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_1227
timestamp 1698431365
transform 1 0 138768 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_1291
timestamp 1698431365
transform 1 0 145936 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_1297
timestamp 1698431365
transform 1 0 146608 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_1361
timestamp 1698431365
transform 1 0 153776 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_1367
timestamp 1698431365
transform 1 0 154448 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_1431
timestamp 1698431365
transform 1 0 161616 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_1437
timestamp 1698431365
transform 1 0 162288 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_1501
timestamp 1698431365
transform 1 0 169456 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_1507
timestamp 1698431365
transform 1 0 170128 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_1571
timestamp 1698431365
transform 1 0 177296 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_1577
timestamp 1698431365
transform 1 0 177968 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_1641
timestamp 1698431365
transform 1 0 185136 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_1647
timestamp 1698431365
transform 1 0 185808 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_1711
timestamp 1698431365
transform 1 0 192976 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_1717
timestamp 1698431365
transform 1 0 193648 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_1781
timestamp 1698431365
transform 1 0 200816 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_1787
timestamp 1698431365
transform 1 0 201488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_1851
timestamp 1698431365
transform 1 0 208656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_1857
timestamp 1698431365
transform 1 0 209328 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_1921
timestamp 1698431365
transform 1 0 216496 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_1927
timestamp 1698431365
transform 1 0 217168 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_1935
timestamp 1698431365
transform 1 0 218064 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_1937
timestamp 1698431365
transform 1 0 218288 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698431365
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_72
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_136
timestamp 1698431365
transform 1 0 16576 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_142
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_206
timestamp 1698431365
transform 1 0 24416 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_212
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_276
timestamp 1698431365
transform 1 0 32256 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_282
timestamp 1698431365
transform 1 0 32928 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_346
timestamp 1698431365
transform 1 0 40096 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_352
timestamp 1698431365
transform 1 0 40768 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_416
timestamp 1698431365
transform 1 0 47936 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_422
timestamp 1698431365
transform 1 0 48608 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_486
timestamp 1698431365
transform 1 0 55776 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_492
timestamp 1698431365
transform 1 0 56448 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_556
timestamp 1698431365
transform 1 0 63616 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_562
timestamp 1698431365
transform 1 0 64288 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_626
timestamp 1698431365
transform 1 0 71456 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_632
timestamp 1698431365
transform 1 0 72128 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_696
timestamp 1698431365
transform 1 0 79296 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_702
timestamp 1698431365
transform 1 0 79968 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_766
timestamp 1698431365
transform 1 0 87136 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_772
timestamp 1698431365
transform 1 0 87808 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_836
timestamp 1698431365
transform 1 0 94976 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_842
timestamp 1698431365
transform 1 0 95648 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_906
timestamp 1698431365
transform 1 0 102816 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_912
timestamp 1698431365
transform 1 0 103488 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_976
timestamp 1698431365
transform 1 0 110656 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_982
timestamp 1698431365
transform 1 0 111328 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_1046
timestamp 1698431365
transform 1 0 118496 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_1052
timestamp 1698431365
transform 1 0 119168 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_1116
timestamp 1698431365
transform 1 0 126336 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_1122
timestamp 1698431365
transform 1 0 127008 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_1186
timestamp 1698431365
transform 1 0 134176 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_1192
timestamp 1698431365
transform 1 0 134848 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_1256
timestamp 1698431365
transform 1 0 142016 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_1262
timestamp 1698431365
transform 1 0 142688 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_1326
timestamp 1698431365
transform 1 0 149856 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_1332
timestamp 1698431365
transform 1 0 150528 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_1396
timestamp 1698431365
transform 1 0 157696 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_1402
timestamp 1698431365
transform 1 0 158368 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_1466
timestamp 1698431365
transform 1 0 165536 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_1472
timestamp 1698431365
transform 1 0 166208 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_1536
timestamp 1698431365
transform 1 0 173376 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_1542
timestamp 1698431365
transform 1 0 174048 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_1606
timestamp 1698431365
transform 1 0 181216 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_1612
timestamp 1698431365
transform 1 0 181888 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_1676
timestamp 1698431365
transform 1 0 189056 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_1682
timestamp 1698431365
transform 1 0 189728 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_1746
timestamp 1698431365
transform 1 0 196896 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_1752
timestamp 1698431365
transform 1 0 197568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_1816
timestamp 1698431365
transform 1 0 204736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_1822
timestamp 1698431365
transform 1 0 205408 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_1886
timestamp 1698431365
transform 1 0 212576 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_1892
timestamp 1698431365
transform 1 0 213248 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_1924
timestamp 1698431365
transform 1 0 216832 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_1932
timestamp 1698431365
transform 1 0 217728 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_1936
timestamp 1698431365
transform 1 0 218176 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698431365
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698431365
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698431365
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_107
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_171
timestamp 1698431365
transform 1 0 20496 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_177
timestamp 1698431365
transform 1 0 21168 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_241
timestamp 1698431365
transform 1 0 28336 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698431365
transform 1 0 29008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698431365
transform 1 0 36176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_317
timestamp 1698431365
transform 1 0 36848 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_381
timestamp 1698431365
transform 1 0 44016 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_387
timestamp 1698431365
transform 1 0 44688 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_451
timestamp 1698431365
transform 1 0 51856 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_457
timestamp 1698431365
transform 1 0 52528 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_521
timestamp 1698431365
transform 1 0 59696 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_527
timestamp 1698431365
transform 1 0 60368 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_591
timestamp 1698431365
transform 1 0 67536 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_597
timestamp 1698431365
transform 1 0 68208 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_661
timestamp 1698431365
transform 1 0 75376 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_667
timestamp 1698431365
transform 1 0 76048 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_731
timestamp 1698431365
transform 1 0 83216 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_737
timestamp 1698431365
transform 1 0 83888 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_801
timestamp 1698431365
transform 1 0 91056 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_807
timestamp 1698431365
transform 1 0 91728 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_871
timestamp 1698431365
transform 1 0 98896 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_877
timestamp 1698431365
transform 1 0 99568 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_941
timestamp 1698431365
transform 1 0 106736 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_947
timestamp 1698431365
transform 1 0 107408 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_1011
timestamp 1698431365
transform 1 0 114576 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_1017
timestamp 1698431365
transform 1 0 115248 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_1081
timestamp 1698431365
transform 1 0 122416 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_1087
timestamp 1698431365
transform 1 0 123088 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_1151
timestamp 1698431365
transform 1 0 130256 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_1157
timestamp 1698431365
transform 1 0 130928 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_1221
timestamp 1698431365
transform 1 0 138096 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_1227
timestamp 1698431365
transform 1 0 138768 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_1291
timestamp 1698431365
transform 1 0 145936 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_1297
timestamp 1698431365
transform 1 0 146608 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_1361
timestamp 1698431365
transform 1 0 153776 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_1367
timestamp 1698431365
transform 1 0 154448 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_1431
timestamp 1698431365
transform 1 0 161616 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_1437
timestamp 1698431365
transform 1 0 162288 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_1501
timestamp 1698431365
transform 1 0 169456 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_1507
timestamp 1698431365
transform 1 0 170128 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_1571
timestamp 1698431365
transform 1 0 177296 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_1577
timestamp 1698431365
transform 1 0 177968 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_1641
timestamp 1698431365
transform 1 0 185136 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_1647
timestamp 1698431365
transform 1 0 185808 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_1711
timestamp 1698431365
transform 1 0 192976 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_1717
timestamp 1698431365
transform 1 0 193648 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_1781
timestamp 1698431365
transform 1 0 200816 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_1787
timestamp 1698431365
transform 1 0 201488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_1851
timestamp 1698431365
transform 1 0 208656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_1857
timestamp 1698431365
transform 1 0 209328 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_1921
timestamp 1698431365
transform 1 0 216496 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_1927
timestamp 1698431365
transform 1 0 217168 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_1935
timestamp 1698431365
transform 1 0 218064 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_1937
timestamp 1698431365
transform 1 0 218288 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698431365
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_72
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_136
timestamp 1698431365
transform 1 0 16576 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_142
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_206
timestamp 1698431365
transform 1 0 24416 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_212
timestamp 1698431365
transform 1 0 25088 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_276
timestamp 1698431365
transform 1 0 32256 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_282
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_346
timestamp 1698431365
transform 1 0 40096 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_352
timestamp 1698431365
transform 1 0 40768 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_416
timestamp 1698431365
transform 1 0 47936 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_422
timestamp 1698431365
transform 1 0 48608 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_486
timestamp 1698431365
transform 1 0 55776 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_492
timestamp 1698431365
transform 1 0 56448 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_556
timestamp 1698431365
transform 1 0 63616 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_562
timestamp 1698431365
transform 1 0 64288 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_626
timestamp 1698431365
transform 1 0 71456 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_632
timestamp 1698431365
transform 1 0 72128 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_696
timestamp 1698431365
transform 1 0 79296 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_702
timestamp 1698431365
transform 1 0 79968 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_766
timestamp 1698431365
transform 1 0 87136 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_772
timestamp 1698431365
transform 1 0 87808 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_836
timestamp 1698431365
transform 1 0 94976 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_842
timestamp 1698431365
transform 1 0 95648 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_906
timestamp 1698431365
transform 1 0 102816 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_912
timestamp 1698431365
transform 1 0 103488 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_976
timestamp 1698431365
transform 1 0 110656 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_982
timestamp 1698431365
transform 1 0 111328 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_1046
timestamp 1698431365
transform 1 0 118496 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_1052
timestamp 1698431365
transform 1 0 119168 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_1116
timestamp 1698431365
transform 1 0 126336 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_1122
timestamp 1698431365
transform 1 0 127008 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_1186
timestamp 1698431365
transform 1 0 134176 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_1192
timestamp 1698431365
transform 1 0 134848 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_1256
timestamp 1698431365
transform 1 0 142016 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_1262
timestamp 1698431365
transform 1 0 142688 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_1326
timestamp 1698431365
transform 1 0 149856 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_1332
timestamp 1698431365
transform 1 0 150528 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_1396
timestamp 1698431365
transform 1 0 157696 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_1402
timestamp 1698431365
transform 1 0 158368 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_1466
timestamp 1698431365
transform 1 0 165536 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_1472
timestamp 1698431365
transform 1 0 166208 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_1536
timestamp 1698431365
transform 1 0 173376 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_1542
timestamp 1698431365
transform 1 0 174048 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_1606
timestamp 1698431365
transform 1 0 181216 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_1612
timestamp 1698431365
transform 1 0 181888 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_1676
timestamp 1698431365
transform 1 0 189056 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_1682
timestamp 1698431365
transform 1 0 189728 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_1746
timestamp 1698431365
transform 1 0 196896 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_1752
timestamp 1698431365
transform 1 0 197568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_1816
timestamp 1698431365
transform 1 0 204736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_1822
timestamp 1698431365
transform 1 0 205408 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_1886
timestamp 1698431365
transform 1 0 212576 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_1892
timestamp 1698431365
transform 1 0 213248 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_1924
timestamp 1698431365
transform 1 0 216832 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_1932
timestamp 1698431365
transform 1 0 217728 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_1936
timestamp 1698431365
transform 1 0 218176 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698431365
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698431365
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698431365
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_107
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_171
timestamp 1698431365
transform 1 0 20496 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_177
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_241
timestamp 1698431365
transform 1 0 28336 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698431365
transform 1 0 36176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_317
timestamp 1698431365
transform 1 0 36848 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_381
timestamp 1698431365
transform 1 0 44016 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_387
timestamp 1698431365
transform 1 0 44688 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_451
timestamp 1698431365
transform 1 0 51856 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_457
timestamp 1698431365
transform 1 0 52528 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_521
timestamp 1698431365
transform 1 0 59696 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_527
timestamp 1698431365
transform 1 0 60368 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_591
timestamp 1698431365
transform 1 0 67536 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_597
timestamp 1698431365
transform 1 0 68208 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_661
timestamp 1698431365
transform 1 0 75376 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_667
timestamp 1698431365
transform 1 0 76048 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_731
timestamp 1698431365
transform 1 0 83216 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_737
timestamp 1698431365
transform 1 0 83888 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_801
timestamp 1698431365
transform 1 0 91056 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_807
timestamp 1698431365
transform 1 0 91728 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_871
timestamp 1698431365
transform 1 0 98896 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_877
timestamp 1698431365
transform 1 0 99568 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_941
timestamp 1698431365
transform 1 0 106736 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_947
timestamp 1698431365
transform 1 0 107408 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_1011
timestamp 1698431365
transform 1 0 114576 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_1017
timestamp 1698431365
transform 1 0 115248 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_1081
timestamp 1698431365
transform 1 0 122416 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_1087
timestamp 1698431365
transform 1 0 123088 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_1151
timestamp 1698431365
transform 1 0 130256 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_1157
timestamp 1698431365
transform 1 0 130928 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_1221
timestamp 1698431365
transform 1 0 138096 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_1227
timestamp 1698431365
transform 1 0 138768 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_1291
timestamp 1698431365
transform 1 0 145936 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_1297
timestamp 1698431365
transform 1 0 146608 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_1361
timestamp 1698431365
transform 1 0 153776 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_1367
timestamp 1698431365
transform 1 0 154448 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_1431
timestamp 1698431365
transform 1 0 161616 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_1437
timestamp 1698431365
transform 1 0 162288 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_1501
timestamp 1698431365
transform 1 0 169456 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_1507
timestamp 1698431365
transform 1 0 170128 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_1571
timestamp 1698431365
transform 1 0 177296 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_1577
timestamp 1698431365
transform 1 0 177968 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_1641
timestamp 1698431365
transform 1 0 185136 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_1647
timestamp 1698431365
transform 1 0 185808 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_1711
timestamp 1698431365
transform 1 0 192976 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_1717
timestamp 1698431365
transform 1 0 193648 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_1781
timestamp 1698431365
transform 1 0 200816 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_1787
timestamp 1698431365
transform 1 0 201488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_1851
timestamp 1698431365
transform 1 0 208656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_1857
timestamp 1698431365
transform 1 0 209328 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_1921
timestamp 1698431365
transform 1 0 216496 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_1927
timestamp 1698431365
transform 1 0 217168 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_1935
timestamp 1698431365
transform 1 0 218064 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_1937
timestamp 1698431365
transform 1 0 218288 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698431365
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_72
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_136
timestamp 1698431365
transform 1 0 16576 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_142
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_206
timestamp 1698431365
transform 1 0 24416 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_212
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_276
timestamp 1698431365
transform 1 0 32256 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_282
timestamp 1698431365
transform 1 0 32928 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_346
timestamp 1698431365
transform 1 0 40096 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_352
timestamp 1698431365
transform 1 0 40768 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_416
timestamp 1698431365
transform 1 0 47936 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_422
timestamp 1698431365
transform 1 0 48608 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_486
timestamp 1698431365
transform 1 0 55776 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_492
timestamp 1698431365
transform 1 0 56448 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_556
timestamp 1698431365
transform 1 0 63616 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_562
timestamp 1698431365
transform 1 0 64288 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_626
timestamp 1698431365
transform 1 0 71456 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_632
timestamp 1698431365
transform 1 0 72128 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_696
timestamp 1698431365
transform 1 0 79296 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_702
timestamp 1698431365
transform 1 0 79968 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_766
timestamp 1698431365
transform 1 0 87136 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_772
timestamp 1698431365
transform 1 0 87808 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_836
timestamp 1698431365
transform 1 0 94976 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_842
timestamp 1698431365
transform 1 0 95648 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_906
timestamp 1698431365
transform 1 0 102816 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_912
timestamp 1698431365
transform 1 0 103488 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_976
timestamp 1698431365
transform 1 0 110656 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_982
timestamp 1698431365
transform 1 0 111328 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_1046
timestamp 1698431365
transform 1 0 118496 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_1052
timestamp 1698431365
transform 1 0 119168 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_1116
timestamp 1698431365
transform 1 0 126336 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_1122
timestamp 1698431365
transform 1 0 127008 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_1186
timestamp 1698431365
transform 1 0 134176 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_1192
timestamp 1698431365
transform 1 0 134848 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_1256
timestamp 1698431365
transform 1 0 142016 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_1262
timestamp 1698431365
transform 1 0 142688 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_1326
timestamp 1698431365
transform 1 0 149856 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_1332
timestamp 1698431365
transform 1 0 150528 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_1396
timestamp 1698431365
transform 1 0 157696 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_1402
timestamp 1698431365
transform 1 0 158368 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_1466
timestamp 1698431365
transform 1 0 165536 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_1472
timestamp 1698431365
transform 1 0 166208 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_1536
timestamp 1698431365
transform 1 0 173376 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_1542
timestamp 1698431365
transform 1 0 174048 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_1606
timestamp 1698431365
transform 1 0 181216 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_1612
timestamp 1698431365
transform 1 0 181888 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_1676
timestamp 1698431365
transform 1 0 189056 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_1682
timestamp 1698431365
transform 1 0 189728 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_1746
timestamp 1698431365
transform 1 0 196896 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_1752
timestamp 1698431365
transform 1 0 197568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_1816
timestamp 1698431365
transform 1 0 204736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_1822
timestamp 1698431365
transform 1 0 205408 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_1886
timestamp 1698431365
transform 1 0 212576 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_1892
timestamp 1698431365
transform 1 0 213248 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_1924
timestamp 1698431365
transform 1 0 216832 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_1932
timestamp 1698431365
transform 1 0 217728 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_1936
timestamp 1698431365
transform 1 0 218176 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698431365
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698431365
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698431365
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_107
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_171
timestamp 1698431365
transform 1 0 20496 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_177
timestamp 1698431365
transform 1 0 21168 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_241
timestamp 1698431365
transform 1 0 28336 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698431365
transform 1 0 29008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698431365
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_317
timestamp 1698431365
transform 1 0 36848 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_381
timestamp 1698431365
transform 1 0 44016 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_387
timestamp 1698431365
transform 1 0 44688 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_451
timestamp 1698431365
transform 1 0 51856 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_457
timestamp 1698431365
transform 1 0 52528 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_521
timestamp 1698431365
transform 1 0 59696 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_527
timestamp 1698431365
transform 1 0 60368 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_591
timestamp 1698431365
transform 1 0 67536 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_597
timestamp 1698431365
transform 1 0 68208 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_661
timestamp 1698431365
transform 1 0 75376 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_667
timestamp 1698431365
transform 1 0 76048 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_731
timestamp 1698431365
transform 1 0 83216 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_737
timestamp 1698431365
transform 1 0 83888 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_801
timestamp 1698431365
transform 1 0 91056 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_807
timestamp 1698431365
transform 1 0 91728 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_871
timestamp 1698431365
transform 1 0 98896 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_877
timestamp 1698431365
transform 1 0 99568 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_941
timestamp 1698431365
transform 1 0 106736 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_947
timestamp 1698431365
transform 1 0 107408 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_1011
timestamp 1698431365
transform 1 0 114576 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_1017
timestamp 1698431365
transform 1 0 115248 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_1081
timestamp 1698431365
transform 1 0 122416 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_1087
timestamp 1698431365
transform 1 0 123088 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_1151
timestamp 1698431365
transform 1 0 130256 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_1157
timestamp 1698431365
transform 1 0 130928 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_1221
timestamp 1698431365
transform 1 0 138096 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_1227
timestamp 1698431365
transform 1 0 138768 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_1291
timestamp 1698431365
transform 1 0 145936 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_1297
timestamp 1698431365
transform 1 0 146608 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_1361
timestamp 1698431365
transform 1 0 153776 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_1367
timestamp 1698431365
transform 1 0 154448 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_1431
timestamp 1698431365
transform 1 0 161616 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_1437
timestamp 1698431365
transform 1 0 162288 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_1501
timestamp 1698431365
transform 1 0 169456 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_1507
timestamp 1698431365
transform 1 0 170128 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_1571
timestamp 1698431365
transform 1 0 177296 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_1577
timestamp 1698431365
transform 1 0 177968 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_1641
timestamp 1698431365
transform 1 0 185136 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_1647
timestamp 1698431365
transform 1 0 185808 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_1711
timestamp 1698431365
transform 1 0 192976 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_1717
timestamp 1698431365
transform 1 0 193648 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_1781
timestamp 1698431365
transform 1 0 200816 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_1787
timestamp 1698431365
transform 1 0 201488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_1851
timestamp 1698431365
transform 1 0 208656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_1857
timestamp 1698431365
transform 1 0 209328 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_1921
timestamp 1698431365
transform 1 0 216496 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_1927
timestamp 1698431365
transform 1 0 217168 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_1935
timestamp 1698431365
transform 1 0 218064 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_1937
timestamp 1698431365
transform 1 0 218288 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698431365
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698431365
transform 1 0 16576 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_142
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_206
timestamp 1698431365
transform 1 0 24416 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698431365
transform 1 0 32256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_346
timestamp 1698431365
transform 1 0 40096 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_352
timestamp 1698431365
transform 1 0 40768 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_416
timestamp 1698431365
transform 1 0 47936 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_422
timestamp 1698431365
transform 1 0 48608 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_486
timestamp 1698431365
transform 1 0 55776 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_492
timestamp 1698431365
transform 1 0 56448 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_556
timestamp 1698431365
transform 1 0 63616 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_562
timestamp 1698431365
transform 1 0 64288 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_626
timestamp 1698431365
transform 1 0 71456 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_632
timestamp 1698431365
transform 1 0 72128 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_696
timestamp 1698431365
transform 1 0 79296 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_702
timestamp 1698431365
transform 1 0 79968 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_766
timestamp 1698431365
transform 1 0 87136 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_772
timestamp 1698431365
transform 1 0 87808 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_836
timestamp 1698431365
transform 1 0 94976 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_842
timestamp 1698431365
transform 1 0 95648 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_906
timestamp 1698431365
transform 1 0 102816 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_912
timestamp 1698431365
transform 1 0 103488 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_976
timestamp 1698431365
transform 1 0 110656 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_982
timestamp 1698431365
transform 1 0 111328 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_1046
timestamp 1698431365
transform 1 0 118496 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_1052
timestamp 1698431365
transform 1 0 119168 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_1116
timestamp 1698431365
transform 1 0 126336 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_1122
timestamp 1698431365
transform 1 0 127008 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_1186
timestamp 1698431365
transform 1 0 134176 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_1192
timestamp 1698431365
transform 1 0 134848 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_1256
timestamp 1698431365
transform 1 0 142016 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_1262
timestamp 1698431365
transform 1 0 142688 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_1326
timestamp 1698431365
transform 1 0 149856 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_1332
timestamp 1698431365
transform 1 0 150528 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_1396
timestamp 1698431365
transform 1 0 157696 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_1402
timestamp 1698431365
transform 1 0 158368 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_1466
timestamp 1698431365
transform 1 0 165536 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_1472
timestamp 1698431365
transform 1 0 166208 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_1536
timestamp 1698431365
transform 1 0 173376 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_1542
timestamp 1698431365
transform 1 0 174048 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_1606
timestamp 1698431365
transform 1 0 181216 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_1612
timestamp 1698431365
transform 1 0 181888 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_1676
timestamp 1698431365
transform 1 0 189056 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_1682
timestamp 1698431365
transform 1 0 189728 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_1746
timestamp 1698431365
transform 1 0 196896 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_1752
timestamp 1698431365
transform 1 0 197568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_1816
timestamp 1698431365
transform 1 0 204736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_1822
timestamp 1698431365
transform 1 0 205408 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_1886
timestamp 1698431365
transform 1 0 212576 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_1892
timestamp 1698431365
transform 1 0 213248 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_1924
timestamp 1698431365
transform 1 0 216832 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_1932
timestamp 1698431365
transform 1 0 217728 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_1936
timestamp 1698431365
transform 1 0 218176 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698431365
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698431365
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698431365
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698431365
transform 1 0 13328 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698431365
transform 1 0 20496 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698431365
transform 1 0 28336 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698431365
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_317
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_381
timestamp 1698431365
transform 1 0 44016 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_387
timestamp 1698431365
transform 1 0 44688 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_451
timestamp 1698431365
transform 1 0 51856 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_457
timestamp 1698431365
transform 1 0 52528 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_521
timestamp 1698431365
transform 1 0 59696 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_527
timestamp 1698431365
transform 1 0 60368 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_591
timestamp 1698431365
transform 1 0 67536 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_597
timestamp 1698431365
transform 1 0 68208 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_661
timestamp 1698431365
transform 1 0 75376 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_667
timestamp 1698431365
transform 1 0 76048 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_731
timestamp 1698431365
transform 1 0 83216 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_737
timestamp 1698431365
transform 1 0 83888 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_801
timestamp 1698431365
transform 1 0 91056 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_807
timestamp 1698431365
transform 1 0 91728 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_871
timestamp 1698431365
transform 1 0 98896 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_877
timestamp 1698431365
transform 1 0 99568 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_941
timestamp 1698431365
transform 1 0 106736 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_947
timestamp 1698431365
transform 1 0 107408 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_1011
timestamp 1698431365
transform 1 0 114576 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_1017
timestamp 1698431365
transform 1 0 115248 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_1081
timestamp 1698431365
transform 1 0 122416 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_1087
timestamp 1698431365
transform 1 0 123088 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_1151
timestamp 1698431365
transform 1 0 130256 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_1157
timestamp 1698431365
transform 1 0 130928 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_1221
timestamp 1698431365
transform 1 0 138096 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_1227
timestamp 1698431365
transform 1 0 138768 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_1291
timestamp 1698431365
transform 1 0 145936 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_1297
timestamp 1698431365
transform 1 0 146608 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_1361
timestamp 1698431365
transform 1 0 153776 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_1367
timestamp 1698431365
transform 1 0 154448 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_1431
timestamp 1698431365
transform 1 0 161616 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_1437
timestamp 1698431365
transform 1 0 162288 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_1501
timestamp 1698431365
transform 1 0 169456 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_1507
timestamp 1698431365
transform 1 0 170128 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_1571
timestamp 1698431365
transform 1 0 177296 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_1577
timestamp 1698431365
transform 1 0 177968 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_1641
timestamp 1698431365
transform 1 0 185136 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_1647
timestamp 1698431365
transform 1 0 185808 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_1711
timestamp 1698431365
transform 1 0 192976 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_1717
timestamp 1698431365
transform 1 0 193648 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_1781
timestamp 1698431365
transform 1 0 200816 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_1787
timestamp 1698431365
transform 1 0 201488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_1851
timestamp 1698431365
transform 1 0 208656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_1857
timestamp 1698431365
transform 1 0 209328 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_1921
timestamp 1698431365
transform 1 0 216496 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_1927
timestamp 1698431365
transform 1 0 217168 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_1935
timestamp 1698431365
transform 1 0 218064 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_1937
timestamp 1698431365
transform 1 0 218288 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698431365
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698431365
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698431365
transform 1 0 17248 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698431365
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698431365
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698431365
transform 1 0 32928 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_346
timestamp 1698431365
transform 1 0 40096 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_352
timestamp 1698431365
transform 1 0 40768 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_416
timestamp 1698431365
transform 1 0 47936 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_422
timestamp 1698431365
transform 1 0 48608 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_486
timestamp 1698431365
transform 1 0 55776 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_492
timestamp 1698431365
transform 1 0 56448 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_556
timestamp 1698431365
transform 1 0 63616 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_562
timestamp 1698431365
transform 1 0 64288 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_626
timestamp 1698431365
transform 1 0 71456 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_632
timestamp 1698431365
transform 1 0 72128 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_696
timestamp 1698431365
transform 1 0 79296 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_702
timestamp 1698431365
transform 1 0 79968 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_766
timestamp 1698431365
transform 1 0 87136 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_772
timestamp 1698431365
transform 1 0 87808 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_836
timestamp 1698431365
transform 1 0 94976 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_842
timestamp 1698431365
transform 1 0 95648 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_858
timestamp 1698431365
transform 1 0 97440 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_860
timestamp 1698431365
transform 1 0 97664 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_890
timestamp 1698431365
transform 1 0 101024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_894
timestamp 1698431365
transform 1 0 101472 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_898
timestamp 1698431365
transform 1 0 101920 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_906
timestamp 1698431365
transform 1 0 102816 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_912
timestamp 1698431365
transform 1 0 103488 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_976
timestamp 1698431365
transform 1 0 110656 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_982
timestamp 1698431365
transform 1 0 111328 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_1046
timestamp 1698431365
transform 1 0 118496 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_1052
timestamp 1698431365
transform 1 0 119168 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_1068
timestamp 1698431365
transform 1 0 120960 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_1101
timestamp 1698431365
transform 1 0 124656 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_1105
timestamp 1698431365
transform 1 0 125104 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_1109
timestamp 1698431365
transform 1 0 125552 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_1117
timestamp 1698431365
transform 1 0 126448 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_1119
timestamp 1698431365
transform 1 0 126672 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_1122
timestamp 1698431365
transform 1 0 127008 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_1154
timestamp 1698431365
transform 1 0 130592 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_1170
timestamp 1698431365
transform 1 0 132384 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_1178
timestamp 1698431365
transform 1 0 133280 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_1182
timestamp 1698431365
transform 1 0 133728 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_1186
timestamp 1698431365
transform 1 0 134176 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_1221
timestamp 1698431365
transform 1 0 138096 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_1253
timestamp 1698431365
transform 1 0 141680 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_1257
timestamp 1698431365
transform 1 0 142128 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_1259
timestamp 1698431365
transform 1 0 142352 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_1262
timestamp 1698431365
transform 1 0 142688 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_1326
timestamp 1698431365
transform 1 0 149856 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_1332
timestamp 1698431365
transform 1 0 150528 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_1396
timestamp 1698431365
transform 1 0 157696 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_1402
timestamp 1698431365
transform 1 0 158368 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_1466
timestamp 1698431365
transform 1 0 165536 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_1472
timestamp 1698431365
transform 1 0 166208 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_1536
timestamp 1698431365
transform 1 0 173376 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_1542
timestamp 1698431365
transform 1 0 174048 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_1606
timestamp 1698431365
transform 1 0 181216 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_1612
timestamp 1698431365
transform 1 0 181888 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_1676
timestamp 1698431365
transform 1 0 189056 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_1682
timestamp 1698431365
transform 1 0 189728 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_1746
timestamp 1698431365
transform 1 0 196896 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_1752
timestamp 1698431365
transform 1 0 197568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_1816
timestamp 1698431365
transform 1 0 204736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_1822
timestamp 1698431365
transform 1 0 205408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_1886
timestamp 1698431365
transform 1 0 212576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_33_1892
timestamp 1698431365
transform 1 0 213248 0 -1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_1924
timestamp 1698431365
transform 1 0 216832 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_1932
timestamp 1698431365
transform 1 0 217728 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_1936
timestamp 1698431365
transform 1 0 218176 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698431365
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698431365
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698431365
transform 1 0 13328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698431365
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698431365
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698431365
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_317
timestamp 1698431365
transform 1 0 36848 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_381
timestamp 1698431365
transform 1 0 44016 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_387
timestamp 1698431365
transform 1 0 44688 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_451
timestamp 1698431365
transform 1 0 51856 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_457
timestamp 1698431365
transform 1 0 52528 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_521
timestamp 1698431365
transform 1 0 59696 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_527
timestamp 1698431365
transform 1 0 60368 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_591
timestamp 1698431365
transform 1 0 67536 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_597
timestamp 1698431365
transform 1 0 68208 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_661
timestamp 1698431365
transform 1 0 75376 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_667
timestamp 1698431365
transform 1 0 76048 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_731
timestamp 1698431365
transform 1 0 83216 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_737
timestamp 1698431365
transform 1 0 83888 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_801
timestamp 1698431365
transform 1 0 91056 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_807
timestamp 1698431365
transform 1 0 91728 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_815
timestamp 1698431365
transform 1 0 92624 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_819
timestamp 1698431365
transform 1 0 93072 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_849
timestamp 1698431365
transform 1 0 96432 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_853
timestamp 1698431365
transform 1 0 96880 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_857
timestamp 1698431365
transform 1 0 97328 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_873
timestamp 1698431365
transform 1 0 99120 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_877
timestamp 1698431365
transform 1 0 99568 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_893
timestamp 1698431365
transform 1 0 101360 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_923
timestamp 1698431365
transform 1 0 104720 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_927
timestamp 1698431365
transform 1 0 105168 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_931
timestamp 1698431365
transform 1 0 105616 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_939
timestamp 1698431365
transform 1 0 106512 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_943
timestamp 1698431365
transform 1 0 106960 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_947
timestamp 1698431365
transform 1 0 107408 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_963
timestamp 1698431365
transform 1 0 109200 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_994
timestamp 1698431365
transform 1 0 112672 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_998
timestamp 1698431365
transform 1 0 113120 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_1002
timestamp 1698431365
transform 1 0 113568 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_1010
timestamp 1698431365
transform 1 0 114464 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_1014
timestamp 1698431365
transform 1 0 114912 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_1017
timestamp 1698431365
transform 1 0 115248 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_1033
timestamp 1698431365
transform 1 0 117040 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_1037
timestamp 1698431365
transform 1 0 117488 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_1069
timestamp 1698431365
transform 1 0 121072 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_1073
timestamp 1698431365
transform 1 0 121520 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_1081
timestamp 1698431365
transform 1 0 122416 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_1087
timestamp 1698431365
transform 1 0 123088 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_1103
timestamp 1698431365
transform 1 0 124880 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_1111
timestamp 1698431365
transform 1 0 125776 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_1142
timestamp 1698431365
transform 1 0 129248 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_1146
timestamp 1698431365
transform 1 0 129696 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_1150
timestamp 1698431365
transform 1 0 130144 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_1154
timestamp 1698431365
transform 1 0 130592 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_1157
timestamp 1698431365
transform 1 0 130928 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_1165
timestamp 1698431365
transform 1 0 131824 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_1169
timestamp 1698431365
transform 1 0 132272 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_1202
timestamp 1698431365
transform 1 0 135968 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_1206
timestamp 1698431365
transform 1 0 136416 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_1222
timestamp 1698431365
transform 1 0 138208 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_1224
timestamp 1698431365
transform 1 0 138432 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_1227
timestamp 1698431365
transform 1 0 138768 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_1291
timestamp 1698431365
transform 1 0 145936 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_1297
timestamp 1698431365
transform 1 0 146608 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_1361
timestamp 1698431365
transform 1 0 153776 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_1367
timestamp 1698431365
transform 1 0 154448 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_1431
timestamp 1698431365
transform 1 0 161616 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_1437
timestamp 1698431365
transform 1 0 162288 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_1501
timestamp 1698431365
transform 1 0 169456 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_1507
timestamp 1698431365
transform 1 0 170128 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_1571
timestamp 1698431365
transform 1 0 177296 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_1577
timestamp 1698431365
transform 1 0 177968 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_1641
timestamp 1698431365
transform 1 0 185136 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_1647
timestamp 1698431365
transform 1 0 185808 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_1711
timestamp 1698431365
transform 1 0 192976 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_1717
timestamp 1698431365
transform 1 0 193648 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_1781
timestamp 1698431365
transform 1 0 200816 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_1787
timestamp 1698431365
transform 1 0 201488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_1851
timestamp 1698431365
transform 1 0 208656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_1857
timestamp 1698431365
transform 1 0 209328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_1921
timestamp 1698431365
transform 1 0 216496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_1927
timestamp 1698431365
transform 1 0 217168 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_1935
timestamp 1698431365
transform 1 0 218064 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_1937
timestamp 1698431365
transform 1 0 218288 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698431365
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698431365
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698431365
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698431365
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698431365
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698431365
transform 1 0 25088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698431365
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_346
timestamp 1698431365
transform 1 0 40096 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_352
timestamp 1698431365
transform 1 0 40768 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_416
timestamp 1698431365
transform 1 0 47936 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_422
timestamp 1698431365
transform 1 0 48608 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_486
timestamp 1698431365
transform 1 0 55776 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_492
timestamp 1698431365
transform 1 0 56448 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_556
timestamp 1698431365
transform 1 0 63616 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_562
timestamp 1698431365
transform 1 0 64288 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_626
timestamp 1698431365
transform 1 0 71456 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_632
timestamp 1698431365
transform 1 0 72128 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_696
timestamp 1698431365
transform 1 0 79296 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_702
timestamp 1698431365
transform 1 0 79968 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_766
timestamp 1698431365
transform 1 0 87136 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_772
timestamp 1698431365
transform 1 0 87808 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_836
timestamp 1698431365
transform 1 0 94976 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_842
timestamp 1698431365
transform 1 0 95648 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_906
timestamp 1698431365
transform 1 0 102816 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_912
timestamp 1698431365
transform 1 0 103488 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_928
timestamp 1698431365
transform 1 0 105280 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_932
timestamp 1698431365
transform 1 0 105728 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_963
timestamp 1698431365
transform 1 0 109200 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_967
timestamp 1698431365
transform 1 0 109648 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_971
timestamp 1698431365
transform 1 0 110096 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_979
timestamp 1698431365
transform 1 0 110992 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_982
timestamp 1698431365
transform 1 0 111328 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_998
timestamp 1698431365
transform 1 0 113120 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_1033
timestamp 1698431365
transform 1 0 117040 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_1037
timestamp 1698431365
transform 1 0 117488 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_1045
timestamp 1698431365
transform 1 0 118384 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_1049
timestamp 1698431365
transform 1 0 118832 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_1052
timestamp 1698431365
transform 1 0 119168 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_1116
timestamp 1698431365
transform 1 0 126336 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_1122
timestamp 1698431365
transform 1 0 127008 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_1186
timestamp 1698431365
transform 1 0 134176 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_1192
timestamp 1698431365
transform 1 0 134848 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_1200
timestamp 1698431365
transform 1 0 135744 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_1204
timestamp 1698431365
transform 1 0 136192 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_1207
timestamp 1698431365
transform 1 0 136528 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_1211
timestamp 1698431365
transform 1 0 136976 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_1242
timestamp 1698431365
transform 1 0 140448 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_1258
timestamp 1698431365
transform 1 0 142240 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_1262
timestamp 1698431365
transform 1 0 142688 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_1326
timestamp 1698431365
transform 1 0 149856 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_1332
timestamp 1698431365
transform 1 0 150528 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_1396
timestamp 1698431365
transform 1 0 157696 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_1402
timestamp 1698431365
transform 1 0 158368 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_1466
timestamp 1698431365
transform 1 0 165536 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_1472
timestamp 1698431365
transform 1 0 166208 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_1536
timestamp 1698431365
transform 1 0 173376 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_1542
timestamp 1698431365
transform 1 0 174048 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_1606
timestamp 1698431365
transform 1 0 181216 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_1612
timestamp 1698431365
transform 1 0 181888 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_1676
timestamp 1698431365
transform 1 0 189056 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_1682
timestamp 1698431365
transform 1 0 189728 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_1746
timestamp 1698431365
transform 1 0 196896 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_1752
timestamp 1698431365
transform 1 0 197568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_1816
timestamp 1698431365
transform 1 0 204736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_1822
timestamp 1698431365
transform 1 0 205408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_1886
timestamp 1698431365
transform 1 0 212576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_1892
timestamp 1698431365
transform 1 0 213248 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_1924
timestamp 1698431365
transform 1 0 216832 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_1932
timestamp 1698431365
transform 1 0 217728 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_1936
timestamp 1698431365
transform 1 0 218176 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698431365
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698431365
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698431365
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698431365
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698431365
transform 1 0 21168 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698431365
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698431365
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_317
timestamp 1698431365
transform 1 0 36848 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_381
timestamp 1698431365
transform 1 0 44016 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_387
timestamp 1698431365
transform 1 0 44688 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_451
timestamp 1698431365
transform 1 0 51856 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_457
timestamp 1698431365
transform 1 0 52528 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_521
timestamp 1698431365
transform 1 0 59696 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_527
timestamp 1698431365
transform 1 0 60368 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_591
timestamp 1698431365
transform 1 0 67536 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_597
timestamp 1698431365
transform 1 0 68208 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_661
timestamp 1698431365
transform 1 0 75376 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_667
timestamp 1698431365
transform 1 0 76048 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_731
timestamp 1698431365
transform 1 0 83216 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_737
timestamp 1698431365
transform 1 0 83888 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_801
timestamp 1698431365
transform 1 0 91056 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_807
timestamp 1698431365
transform 1 0 91728 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_871
timestamp 1698431365
transform 1 0 98896 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_877
timestamp 1698431365
transform 1 0 99568 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_941
timestamp 1698431365
transform 1 0 106736 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_947
timestamp 1698431365
transform 1 0 107408 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_1011
timestamp 1698431365
transform 1 0 114576 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_1017
timestamp 1698431365
transform 1 0 115248 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_1081
timestamp 1698431365
transform 1 0 122416 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_1087
timestamp 1698431365
transform 1 0 123088 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_1151
timestamp 1698431365
transform 1 0 130256 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_1157
timestamp 1698431365
transform 1 0 130928 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_1221
timestamp 1698431365
transform 1 0 138096 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_1227
timestamp 1698431365
transform 1 0 138768 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_1291
timestamp 1698431365
transform 1 0 145936 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_1297
timestamp 1698431365
transform 1 0 146608 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_1361
timestamp 1698431365
transform 1 0 153776 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_1367
timestamp 1698431365
transform 1 0 154448 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_1431
timestamp 1698431365
transform 1 0 161616 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_1437
timestamp 1698431365
transform 1 0 162288 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_1501
timestamp 1698431365
transform 1 0 169456 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_1507
timestamp 1698431365
transform 1 0 170128 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_1571
timestamp 1698431365
transform 1 0 177296 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_1577
timestamp 1698431365
transform 1 0 177968 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_1641
timestamp 1698431365
transform 1 0 185136 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_1647
timestamp 1698431365
transform 1 0 185808 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_1711
timestamp 1698431365
transform 1 0 192976 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_1717
timestamp 1698431365
transform 1 0 193648 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_1781
timestamp 1698431365
transform 1 0 200816 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_1787
timestamp 1698431365
transform 1 0 201488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_1851
timestamp 1698431365
transform 1 0 208656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_1857
timestamp 1698431365
transform 1 0 209328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_1921
timestamp 1698431365
transform 1 0 216496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_1927
timestamp 1698431365
transform 1 0 217168 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_1935
timestamp 1698431365
transform 1 0 218064 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_1937
timestamp 1698431365
transform 1 0 218288 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698431365
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698431365
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698431365
transform 1 0 17248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698431365
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698431365
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698431365
transform 1 0 32928 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_346
timestamp 1698431365
transform 1 0 40096 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_352
timestamp 1698431365
transform 1 0 40768 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_416
timestamp 1698431365
transform 1 0 47936 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_422
timestamp 1698431365
transform 1 0 48608 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_486
timestamp 1698431365
transform 1 0 55776 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_492
timestamp 1698431365
transform 1 0 56448 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_556
timestamp 1698431365
transform 1 0 63616 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_562
timestamp 1698431365
transform 1 0 64288 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_626
timestamp 1698431365
transform 1 0 71456 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_632
timestamp 1698431365
transform 1 0 72128 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_696
timestamp 1698431365
transform 1 0 79296 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_702
timestamp 1698431365
transform 1 0 79968 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_766
timestamp 1698431365
transform 1 0 87136 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_772
timestamp 1698431365
transform 1 0 87808 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_836
timestamp 1698431365
transform 1 0 94976 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_842
timestamp 1698431365
transform 1 0 95648 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_906
timestamp 1698431365
transform 1 0 102816 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_912
timestamp 1698431365
transform 1 0 103488 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_976
timestamp 1698431365
transform 1 0 110656 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_1032
timestamp 1698431365
transform 1 0 116928 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_1036
timestamp 1698431365
transform 1 0 117376 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_1044
timestamp 1698431365
transform 1 0 118272 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_1048
timestamp 1698431365
transform 1 0 118720 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_1052
timestamp 1698431365
transform 1 0 119168 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_1116
timestamp 1698431365
transform 1 0 126336 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_1122
timestamp 1698431365
transform 1 0 127008 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_1186
timestamp 1698431365
transform 1 0 134176 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_1192
timestamp 1698431365
transform 1 0 134848 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_1256
timestamp 1698431365
transform 1 0 142016 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_1262
timestamp 1698431365
transform 1 0 142688 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_1326
timestamp 1698431365
transform 1 0 149856 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_1332
timestamp 1698431365
transform 1 0 150528 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_1396
timestamp 1698431365
transform 1 0 157696 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_1402
timestamp 1698431365
transform 1 0 158368 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_1466
timestamp 1698431365
transform 1 0 165536 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_1472
timestamp 1698431365
transform 1 0 166208 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_1536
timestamp 1698431365
transform 1 0 173376 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_1542
timestamp 1698431365
transform 1 0 174048 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_1606
timestamp 1698431365
transform 1 0 181216 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_1612
timestamp 1698431365
transform 1 0 181888 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_1676
timestamp 1698431365
transform 1 0 189056 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_1682
timestamp 1698431365
transform 1 0 189728 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_1746
timestamp 1698431365
transform 1 0 196896 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_1752
timestamp 1698431365
transform 1 0 197568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_1816
timestamp 1698431365
transform 1 0 204736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_1822
timestamp 1698431365
transform 1 0 205408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_1886
timestamp 1698431365
transform 1 0 212576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_1892
timestamp 1698431365
transform 1 0 213248 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_1924
timestamp 1698431365
transform 1 0 216832 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_1932
timestamp 1698431365
transform 1 0 217728 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_1936
timestamp 1698431365
transform 1 0 218176 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698431365
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698431365
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698431365
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698431365
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698431365
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698431365
transform 1 0 29008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698431365
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_317
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_381
timestamp 1698431365
transform 1 0 44016 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_387
timestamp 1698431365
transform 1 0 44688 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_451
timestamp 1698431365
transform 1 0 51856 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_457
timestamp 1698431365
transform 1 0 52528 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_521
timestamp 1698431365
transform 1 0 59696 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_527
timestamp 1698431365
transform 1 0 60368 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_591
timestamp 1698431365
transform 1 0 67536 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_597
timestamp 1698431365
transform 1 0 68208 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_661
timestamp 1698431365
transform 1 0 75376 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_667
timestamp 1698431365
transform 1 0 76048 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_731
timestamp 1698431365
transform 1 0 83216 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_737
timestamp 1698431365
transform 1 0 83888 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_801
timestamp 1698431365
transform 1 0 91056 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_807
timestamp 1698431365
transform 1 0 91728 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_871
timestamp 1698431365
transform 1 0 98896 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_877
timestamp 1698431365
transform 1 0 99568 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_941
timestamp 1698431365
transform 1 0 106736 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_947
timestamp 1698431365
transform 1 0 107408 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_1011
timestamp 1698431365
transform 1 0 114576 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_1017
timestamp 1698431365
transform 1 0 115248 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_1081
timestamp 1698431365
transform 1 0 122416 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_1087
timestamp 1698431365
transform 1 0 123088 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_1151
timestamp 1698431365
transform 1 0 130256 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_1157
timestamp 1698431365
transform 1 0 130928 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_1221
timestamp 1698431365
transform 1 0 138096 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_1227
timestamp 1698431365
transform 1 0 138768 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_1291
timestamp 1698431365
transform 1 0 145936 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_1297
timestamp 1698431365
transform 1 0 146608 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_1361
timestamp 1698431365
transform 1 0 153776 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_1367
timestamp 1698431365
transform 1 0 154448 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_1431
timestamp 1698431365
transform 1 0 161616 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_1437
timestamp 1698431365
transform 1 0 162288 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_1501
timestamp 1698431365
transform 1 0 169456 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_1507
timestamp 1698431365
transform 1 0 170128 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_1571
timestamp 1698431365
transform 1 0 177296 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_1577
timestamp 1698431365
transform 1 0 177968 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_1641
timestamp 1698431365
transform 1 0 185136 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_1647
timestamp 1698431365
transform 1 0 185808 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_1711
timestamp 1698431365
transform 1 0 192976 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_1717
timestamp 1698431365
transform 1 0 193648 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_1781
timestamp 1698431365
transform 1 0 200816 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_1787
timestamp 1698431365
transform 1 0 201488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_1851
timestamp 1698431365
transform 1 0 208656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_1857
timestamp 1698431365
transform 1 0 209328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_1921
timestamp 1698431365
transform 1 0 216496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_1927
timestamp 1698431365
transform 1 0 217168 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_1935
timestamp 1698431365
transform 1 0 218064 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_1937
timestamp 1698431365
transform 1 0 218288 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698431365
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698431365
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698431365
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698431365
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698431365
transform 1 0 32928 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_346
timestamp 1698431365
transform 1 0 40096 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_352
timestamp 1698431365
transform 1 0 40768 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_416
timestamp 1698431365
transform 1 0 47936 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_422
timestamp 1698431365
transform 1 0 48608 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_486
timestamp 1698431365
transform 1 0 55776 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_492
timestamp 1698431365
transform 1 0 56448 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_556
timestamp 1698431365
transform 1 0 63616 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_562
timestamp 1698431365
transform 1 0 64288 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_626
timestamp 1698431365
transform 1 0 71456 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_632
timestamp 1698431365
transform 1 0 72128 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_696
timestamp 1698431365
transform 1 0 79296 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_702
timestamp 1698431365
transform 1 0 79968 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_766
timestamp 1698431365
transform 1 0 87136 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_772
timestamp 1698431365
transform 1 0 87808 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_836
timestamp 1698431365
transform 1 0 94976 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_842
timestamp 1698431365
transform 1 0 95648 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_906
timestamp 1698431365
transform 1 0 102816 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_912
timestamp 1698431365
transform 1 0 103488 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_976
timestamp 1698431365
transform 1 0 110656 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_982
timestamp 1698431365
transform 1 0 111328 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_1046
timestamp 1698431365
transform 1 0 118496 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_1052
timestamp 1698431365
transform 1 0 119168 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_1116
timestamp 1698431365
transform 1 0 126336 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_1122
timestamp 1698431365
transform 1 0 127008 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_1186
timestamp 1698431365
transform 1 0 134176 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_1192
timestamp 1698431365
transform 1 0 134848 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_1256
timestamp 1698431365
transform 1 0 142016 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_1262
timestamp 1698431365
transform 1 0 142688 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_1326
timestamp 1698431365
transform 1 0 149856 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_1332
timestamp 1698431365
transform 1 0 150528 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_1396
timestamp 1698431365
transform 1 0 157696 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_1402
timestamp 1698431365
transform 1 0 158368 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_1466
timestamp 1698431365
transform 1 0 165536 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_1472
timestamp 1698431365
transform 1 0 166208 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_1536
timestamp 1698431365
transform 1 0 173376 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_1542
timestamp 1698431365
transform 1 0 174048 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_1606
timestamp 1698431365
transform 1 0 181216 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_1612
timestamp 1698431365
transform 1 0 181888 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_1676
timestamp 1698431365
transform 1 0 189056 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_1682
timestamp 1698431365
transform 1 0 189728 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_1746
timestamp 1698431365
transform 1 0 196896 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_1752
timestamp 1698431365
transform 1 0 197568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_1816
timestamp 1698431365
transform 1 0 204736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_1822
timestamp 1698431365
transform 1 0 205408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_1886
timestamp 1698431365
transform 1 0 212576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_1892
timestamp 1698431365
transform 1 0 213248 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_1924
timestamp 1698431365
transform 1 0 216832 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_1932
timestamp 1698431365
transform 1 0 217728 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_1936
timestamp 1698431365
transform 1 0 218176 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698431365
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698431365
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698431365
transform 1 0 13328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698431365
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698431365
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698431365
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_317
timestamp 1698431365
transform 1 0 36848 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_381
timestamp 1698431365
transform 1 0 44016 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_387
timestamp 1698431365
transform 1 0 44688 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_451
timestamp 1698431365
transform 1 0 51856 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_457
timestamp 1698431365
transform 1 0 52528 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_521
timestamp 1698431365
transform 1 0 59696 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_527
timestamp 1698431365
transform 1 0 60368 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_591
timestamp 1698431365
transform 1 0 67536 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_597
timestamp 1698431365
transform 1 0 68208 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_661
timestamp 1698431365
transform 1 0 75376 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_667
timestamp 1698431365
transform 1 0 76048 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_731
timestamp 1698431365
transform 1 0 83216 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_737
timestamp 1698431365
transform 1 0 83888 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_801
timestamp 1698431365
transform 1 0 91056 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_807
timestamp 1698431365
transform 1 0 91728 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_871
timestamp 1698431365
transform 1 0 98896 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_877
timestamp 1698431365
transform 1 0 99568 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_941
timestamp 1698431365
transform 1 0 106736 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_947
timestamp 1698431365
transform 1 0 107408 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_1011
timestamp 1698431365
transform 1 0 114576 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_1017
timestamp 1698431365
transform 1 0 115248 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_1081
timestamp 1698431365
transform 1 0 122416 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_1087
timestamp 1698431365
transform 1 0 123088 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_1151
timestamp 1698431365
transform 1 0 130256 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_1157
timestamp 1698431365
transform 1 0 130928 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_1221
timestamp 1698431365
transform 1 0 138096 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_1227
timestamp 1698431365
transform 1 0 138768 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_1291
timestamp 1698431365
transform 1 0 145936 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_1297
timestamp 1698431365
transform 1 0 146608 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_1361
timestamp 1698431365
transform 1 0 153776 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_1367
timestamp 1698431365
transform 1 0 154448 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_1431
timestamp 1698431365
transform 1 0 161616 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_1437
timestamp 1698431365
transform 1 0 162288 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_1501
timestamp 1698431365
transform 1 0 169456 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_1507
timestamp 1698431365
transform 1 0 170128 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_1571
timestamp 1698431365
transform 1 0 177296 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_1577
timestamp 1698431365
transform 1 0 177968 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_1641
timestamp 1698431365
transform 1 0 185136 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_1647
timestamp 1698431365
transform 1 0 185808 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_1711
timestamp 1698431365
transform 1 0 192976 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_1717
timestamp 1698431365
transform 1 0 193648 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_1781
timestamp 1698431365
transform 1 0 200816 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_1787
timestamp 1698431365
transform 1 0 201488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_1851
timestamp 1698431365
transform 1 0 208656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_1857
timestamp 1698431365
transform 1 0 209328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_1921
timestamp 1698431365
transform 1 0 216496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_1927
timestamp 1698431365
transform 1 0 217168 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_1935
timestamp 1698431365
transform 1 0 218064 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_1937
timestamp 1698431365
transform 1 0 218288 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698431365
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698431365
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698431365
transform 1 0 17248 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698431365
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698431365
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698431365
transform 1 0 32928 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_346
timestamp 1698431365
transform 1 0 40096 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_352
timestamp 1698431365
transform 1 0 40768 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_416
timestamp 1698431365
transform 1 0 47936 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_422
timestamp 1698431365
transform 1 0 48608 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_486
timestamp 1698431365
transform 1 0 55776 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_492
timestamp 1698431365
transform 1 0 56448 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_556
timestamp 1698431365
transform 1 0 63616 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_562
timestamp 1698431365
transform 1 0 64288 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_626
timestamp 1698431365
transform 1 0 71456 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_632
timestamp 1698431365
transform 1 0 72128 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_696
timestamp 1698431365
transform 1 0 79296 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_702
timestamp 1698431365
transform 1 0 79968 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_766
timestamp 1698431365
transform 1 0 87136 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_772
timestamp 1698431365
transform 1 0 87808 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_836
timestamp 1698431365
transform 1 0 94976 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_842
timestamp 1698431365
transform 1 0 95648 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_906
timestamp 1698431365
transform 1 0 102816 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_912
timestamp 1698431365
transform 1 0 103488 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_976
timestamp 1698431365
transform 1 0 110656 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_982
timestamp 1698431365
transform 1 0 111328 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_1046
timestamp 1698431365
transform 1 0 118496 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_1052
timestamp 1698431365
transform 1 0 119168 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_1116
timestamp 1698431365
transform 1 0 126336 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_1122
timestamp 1698431365
transform 1 0 127008 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_1186
timestamp 1698431365
transform 1 0 134176 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_1192
timestamp 1698431365
transform 1 0 134848 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_1256
timestamp 1698431365
transform 1 0 142016 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_1262
timestamp 1698431365
transform 1 0 142688 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_1326
timestamp 1698431365
transform 1 0 149856 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_1332
timestamp 1698431365
transform 1 0 150528 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_1396
timestamp 1698431365
transform 1 0 157696 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_1402
timestamp 1698431365
transform 1 0 158368 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_1466
timestamp 1698431365
transform 1 0 165536 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_1472
timestamp 1698431365
transform 1 0 166208 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_1536
timestamp 1698431365
transform 1 0 173376 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_1542
timestamp 1698431365
transform 1 0 174048 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_1606
timestamp 1698431365
transform 1 0 181216 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_1612
timestamp 1698431365
transform 1 0 181888 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_1676
timestamp 1698431365
transform 1 0 189056 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_1682
timestamp 1698431365
transform 1 0 189728 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_1746
timestamp 1698431365
transform 1 0 196896 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_1752
timestamp 1698431365
transform 1 0 197568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_1816
timestamp 1698431365
transform 1 0 204736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_1822
timestamp 1698431365
transform 1 0 205408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_1886
timestamp 1698431365
transform 1 0 212576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_1892
timestamp 1698431365
transform 1 0 213248 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_1924
timestamp 1698431365
transform 1 0 216832 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_1932
timestamp 1698431365
transform 1 0 217728 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_1936
timestamp 1698431365
transform 1 0 218176 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698431365
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698431365
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698431365
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698431365
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698431365
transform 1 0 13328 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698431365
transform 1 0 20496 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698431365
transform 1 0 21168 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698431365
transform 1 0 28336 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698431365
transform 1 0 29008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698431365
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_317
timestamp 1698431365
transform 1 0 36848 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_381
timestamp 1698431365
transform 1 0 44016 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_387
timestamp 1698431365
transform 1 0 44688 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_451
timestamp 1698431365
transform 1 0 51856 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_457
timestamp 1698431365
transform 1 0 52528 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_521
timestamp 1698431365
transform 1 0 59696 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_527
timestamp 1698431365
transform 1 0 60368 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_591
timestamp 1698431365
transform 1 0 67536 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_597
timestamp 1698431365
transform 1 0 68208 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_661
timestamp 1698431365
transform 1 0 75376 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_667
timestamp 1698431365
transform 1 0 76048 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_731
timestamp 1698431365
transform 1 0 83216 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_737
timestamp 1698431365
transform 1 0 83888 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_801
timestamp 1698431365
transform 1 0 91056 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_807
timestamp 1698431365
transform 1 0 91728 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_871
timestamp 1698431365
transform 1 0 98896 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_877
timestamp 1698431365
transform 1 0 99568 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_941
timestamp 1698431365
transform 1 0 106736 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_947
timestamp 1698431365
transform 1 0 107408 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_1011
timestamp 1698431365
transform 1 0 114576 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_1017
timestamp 1698431365
transform 1 0 115248 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_1081
timestamp 1698431365
transform 1 0 122416 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_1087
timestamp 1698431365
transform 1 0 123088 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_1151
timestamp 1698431365
transform 1 0 130256 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_1207
timestamp 1698431365
transform 1 0 136528 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_1223
timestamp 1698431365
transform 1 0 138320 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_1227
timestamp 1698431365
transform 1 0 138768 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_1291
timestamp 1698431365
transform 1 0 145936 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_1297
timestamp 1698431365
transform 1 0 146608 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_1361
timestamp 1698431365
transform 1 0 153776 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_1367
timestamp 1698431365
transform 1 0 154448 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_1431
timestamp 1698431365
transform 1 0 161616 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_1437
timestamp 1698431365
transform 1 0 162288 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_1501
timestamp 1698431365
transform 1 0 169456 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_1507
timestamp 1698431365
transform 1 0 170128 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_1571
timestamp 1698431365
transform 1 0 177296 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_1577
timestamp 1698431365
transform 1 0 177968 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_1641
timestamp 1698431365
transform 1 0 185136 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_1647
timestamp 1698431365
transform 1 0 185808 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_1711
timestamp 1698431365
transform 1 0 192976 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_1717
timestamp 1698431365
transform 1 0 193648 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_1781
timestamp 1698431365
transform 1 0 200816 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_1787
timestamp 1698431365
transform 1 0 201488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_1851
timestamp 1698431365
transform 1 0 208656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_1857
timestamp 1698431365
transform 1 0 209328 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_1921
timestamp 1698431365
transform 1 0 216496 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_1927
timestamp 1698431365
transform 1 0 217168 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_1935
timestamp 1698431365
transform 1 0 218064 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_1937
timestamp 1698431365
transform 1 0 218288 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698431365
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698431365
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698431365
transform 1 0 9408 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698431365
transform 1 0 16576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_142
timestamp 1698431365
transform 1 0 17248 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_206
timestamp 1698431365
transform 1 0 24416 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_212
timestamp 1698431365
transform 1 0 25088 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_276
timestamp 1698431365
transform 1 0 32256 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698431365
transform 1 0 32928 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_346
timestamp 1698431365
transform 1 0 40096 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_352
timestamp 1698431365
transform 1 0 40768 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_416
timestamp 1698431365
transform 1 0 47936 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_422
timestamp 1698431365
transform 1 0 48608 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_486
timestamp 1698431365
transform 1 0 55776 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_492
timestamp 1698431365
transform 1 0 56448 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_556
timestamp 1698431365
transform 1 0 63616 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_562
timestamp 1698431365
transform 1 0 64288 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_626
timestamp 1698431365
transform 1 0 71456 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_632
timestamp 1698431365
transform 1 0 72128 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_696
timestamp 1698431365
transform 1 0 79296 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_702
timestamp 1698431365
transform 1 0 79968 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_766
timestamp 1698431365
transform 1 0 87136 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_772
timestamp 1698431365
transform 1 0 87808 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_836
timestamp 1698431365
transform 1 0 94976 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_842
timestamp 1698431365
transform 1 0 95648 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_906
timestamp 1698431365
transform 1 0 102816 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_912
timestamp 1698431365
transform 1 0 103488 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_976
timestamp 1698431365
transform 1 0 110656 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_982
timestamp 1698431365
transform 1 0 111328 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_1046
timestamp 1698431365
transform 1 0 118496 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_1102
timestamp 1698431365
transform 1 0 124768 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_1118
timestamp 1698431365
transform 1 0 126560 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_1122
timestamp 1698431365
transform 1 0 127008 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_1186
timestamp 1698431365
transform 1 0 134176 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_1192
timestamp 1698431365
transform 1 0 134848 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_1256
timestamp 1698431365
transform 1 0 142016 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_1262
timestamp 1698431365
transform 1 0 142688 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_1326
timestamp 1698431365
transform 1 0 149856 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_1332
timestamp 1698431365
transform 1 0 150528 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_1396
timestamp 1698431365
transform 1 0 157696 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_1402
timestamp 1698431365
transform 1 0 158368 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_1466
timestamp 1698431365
transform 1 0 165536 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_1472
timestamp 1698431365
transform 1 0 166208 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_1536
timestamp 1698431365
transform 1 0 173376 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_1542
timestamp 1698431365
transform 1 0 174048 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_1606
timestamp 1698431365
transform 1 0 181216 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_1612
timestamp 1698431365
transform 1 0 181888 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_1676
timestamp 1698431365
transform 1 0 189056 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_1682
timestamp 1698431365
transform 1 0 189728 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_1746
timestamp 1698431365
transform 1 0 196896 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_1752
timestamp 1698431365
transform 1 0 197568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_1816
timestamp 1698431365
transform 1 0 204736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_1822
timestamp 1698431365
transform 1 0 205408 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_1886
timestamp 1698431365
transform 1 0 212576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_1892
timestamp 1698431365
transform 1 0 213248 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_1924
timestamp 1698431365
transform 1 0 216832 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_1932
timestamp 1698431365
transform 1 0 217728 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_1936
timestamp 1698431365
transform 1 0 218176 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698431365
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_34
timestamp 1698431365
transform 1 0 5152 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_37
timestamp 1698431365
transform 1 0 5488 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_101
timestamp 1698431365
transform 1 0 12656 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_107
timestamp 1698431365
transform 1 0 13328 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_171
timestamp 1698431365
transform 1 0 20496 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_177
timestamp 1698431365
transform 1 0 21168 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_241
timestamp 1698431365
transform 1 0 28336 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_247
timestamp 1698431365
transform 1 0 29008 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_311
timestamp 1698431365
transform 1 0 36176 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_317
timestamp 1698431365
transform 1 0 36848 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_381
timestamp 1698431365
transform 1 0 44016 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_387
timestamp 1698431365
transform 1 0 44688 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_451
timestamp 1698431365
transform 1 0 51856 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_457
timestamp 1698431365
transform 1 0 52528 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_521
timestamp 1698431365
transform 1 0 59696 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_527
timestamp 1698431365
transform 1 0 60368 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_591
timestamp 1698431365
transform 1 0 67536 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_597
timestamp 1698431365
transform 1 0 68208 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_661
timestamp 1698431365
transform 1 0 75376 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_667
timestamp 1698431365
transform 1 0 76048 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_731
timestamp 1698431365
transform 1 0 83216 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_737
timestamp 1698431365
transform 1 0 83888 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_801
timestamp 1698431365
transform 1 0 91056 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_807
timestamp 1698431365
transform 1 0 91728 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_871
timestamp 1698431365
transform 1 0 98896 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_877
timestamp 1698431365
transform 1 0 99568 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_941
timestamp 1698431365
transform 1 0 106736 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_947
timestamp 1698431365
transform 1 0 107408 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_1011
timestamp 1698431365
transform 1 0 114576 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_1017
timestamp 1698431365
transform 1 0 115248 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_1081
timestamp 1698431365
transform 1 0 122416 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_1087
timestamp 1698431365
transform 1 0 123088 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_1151
timestamp 1698431365
transform 1 0 130256 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_1157
timestamp 1698431365
transform 1 0 130928 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_1221
timestamp 1698431365
transform 1 0 138096 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_1227
timestamp 1698431365
transform 1 0 138768 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_1291
timestamp 1698431365
transform 1 0 145936 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_1297
timestamp 1698431365
transform 1 0 146608 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_1361
timestamp 1698431365
transform 1 0 153776 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_1367
timestamp 1698431365
transform 1 0 154448 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_1431
timestamp 1698431365
transform 1 0 161616 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_1437
timestamp 1698431365
transform 1 0 162288 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_1501
timestamp 1698431365
transform 1 0 169456 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_1507
timestamp 1698431365
transform 1 0 170128 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_1571
timestamp 1698431365
transform 1 0 177296 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_1577
timestamp 1698431365
transform 1 0 177968 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_1641
timestamp 1698431365
transform 1 0 185136 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_1647
timestamp 1698431365
transform 1 0 185808 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_1711
timestamp 1698431365
transform 1 0 192976 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_1717
timestamp 1698431365
transform 1 0 193648 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_1781
timestamp 1698431365
transform 1 0 200816 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_1787
timestamp 1698431365
transform 1 0 201488 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_1851
timestamp 1698431365
transform 1 0 208656 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_44_1857
timestamp 1698431365
transform 1 0 209328 0 1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_1921
timestamp 1698431365
transform 1 0 216496 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_1927
timestamp 1698431365
transform 1 0 217168 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_1935
timestamp 1698431365
transform 1 0 218064 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_1937
timestamp 1698431365
transform 1 0 218288 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_2
timestamp 1698431365
transform 1 0 1568 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_66
timestamp 1698431365
transform 1 0 8736 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_72
timestamp 1698431365
transform 1 0 9408 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_136
timestamp 1698431365
transform 1 0 16576 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_142
timestamp 1698431365
transform 1 0 17248 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_206
timestamp 1698431365
transform 1 0 24416 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_212
timestamp 1698431365
transform 1 0 25088 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_276
timestamp 1698431365
transform 1 0 32256 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_282
timestamp 1698431365
transform 1 0 32928 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_346
timestamp 1698431365
transform 1 0 40096 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_352
timestamp 1698431365
transform 1 0 40768 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_416
timestamp 1698431365
transform 1 0 47936 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_422
timestamp 1698431365
transform 1 0 48608 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_486
timestamp 1698431365
transform 1 0 55776 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_492
timestamp 1698431365
transform 1 0 56448 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_556
timestamp 1698431365
transform 1 0 63616 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_562
timestamp 1698431365
transform 1 0 64288 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_626
timestamp 1698431365
transform 1 0 71456 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_632
timestamp 1698431365
transform 1 0 72128 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_696
timestamp 1698431365
transform 1 0 79296 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_702
timestamp 1698431365
transform 1 0 79968 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_766
timestamp 1698431365
transform 1 0 87136 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_772
timestamp 1698431365
transform 1 0 87808 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_836
timestamp 1698431365
transform 1 0 94976 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_842
timestamp 1698431365
transform 1 0 95648 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_906
timestamp 1698431365
transform 1 0 102816 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_912
timestamp 1698431365
transform 1 0 103488 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_976
timestamp 1698431365
transform 1 0 110656 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_982
timestamp 1698431365
transform 1 0 111328 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_1046
timestamp 1698431365
transform 1 0 118496 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_1052
timestamp 1698431365
transform 1 0 119168 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_1116
timestamp 1698431365
transform 1 0 126336 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_1122
timestamp 1698431365
transform 1 0 127008 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_1186
timestamp 1698431365
transform 1 0 134176 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_1192
timestamp 1698431365
transform 1 0 134848 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_1256
timestamp 1698431365
transform 1 0 142016 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_1262
timestamp 1698431365
transform 1 0 142688 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_1326
timestamp 1698431365
transform 1 0 149856 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_1332
timestamp 1698431365
transform 1 0 150528 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_1396
timestamp 1698431365
transform 1 0 157696 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_1402
timestamp 1698431365
transform 1 0 158368 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_1466
timestamp 1698431365
transform 1 0 165536 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_1472
timestamp 1698431365
transform 1 0 166208 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_1536
timestamp 1698431365
transform 1 0 173376 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_1542
timestamp 1698431365
transform 1 0 174048 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_1606
timestamp 1698431365
transform 1 0 181216 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_1612
timestamp 1698431365
transform 1 0 181888 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_1676
timestamp 1698431365
transform 1 0 189056 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_1682
timestamp 1698431365
transform 1 0 189728 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_1746
timestamp 1698431365
transform 1 0 196896 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_1752
timestamp 1698431365
transform 1 0 197568 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_1816
timestamp 1698431365
transform 1 0 204736 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_45_1822
timestamp 1698431365
transform 1 0 205408 0 -1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_1886
timestamp 1698431365
transform 1 0 212576 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_1892
timestamp 1698431365
transform 1 0 213248 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_1924
timestamp 1698431365
transform 1 0 216832 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_1932
timestamp 1698431365
transform 1 0 217728 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_1936
timestamp 1698431365
transform 1 0 218176 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_2
timestamp 1698431365
transform 1 0 1568 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_34
timestamp 1698431365
transform 1 0 5152 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_37
timestamp 1698431365
transform 1 0 5488 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_101
timestamp 1698431365
transform 1 0 12656 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_107
timestamp 1698431365
transform 1 0 13328 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_171
timestamp 1698431365
transform 1 0 20496 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_177
timestamp 1698431365
transform 1 0 21168 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_241
timestamp 1698431365
transform 1 0 28336 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_247
timestamp 1698431365
transform 1 0 29008 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_311
timestamp 1698431365
transform 1 0 36176 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_317
timestamp 1698431365
transform 1 0 36848 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_381
timestamp 1698431365
transform 1 0 44016 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_387
timestamp 1698431365
transform 1 0 44688 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_451
timestamp 1698431365
transform 1 0 51856 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_457
timestamp 1698431365
transform 1 0 52528 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_521
timestamp 1698431365
transform 1 0 59696 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_527
timestamp 1698431365
transform 1 0 60368 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_591
timestamp 1698431365
transform 1 0 67536 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_597
timestamp 1698431365
transform 1 0 68208 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_661
timestamp 1698431365
transform 1 0 75376 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_667
timestamp 1698431365
transform 1 0 76048 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_731
timestamp 1698431365
transform 1 0 83216 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_737
timestamp 1698431365
transform 1 0 83888 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_801
timestamp 1698431365
transform 1 0 91056 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_807
timestamp 1698431365
transform 1 0 91728 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_871
timestamp 1698431365
transform 1 0 98896 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_877
timestamp 1698431365
transform 1 0 99568 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_941
timestamp 1698431365
transform 1 0 106736 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_947
timestamp 1698431365
transform 1 0 107408 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_1011
timestamp 1698431365
transform 1 0 114576 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_1017
timestamp 1698431365
transform 1 0 115248 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_1081
timestamp 1698431365
transform 1 0 122416 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_1087
timestamp 1698431365
transform 1 0 123088 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_1151
timestamp 1698431365
transform 1 0 130256 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_1157
timestamp 1698431365
transform 1 0 130928 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_1221
timestamp 1698431365
transform 1 0 138096 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_1227
timestamp 1698431365
transform 1 0 138768 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_1291
timestamp 1698431365
transform 1 0 145936 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_1297
timestamp 1698431365
transform 1 0 146608 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_1361
timestamp 1698431365
transform 1 0 153776 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_1367
timestamp 1698431365
transform 1 0 154448 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_1431
timestamp 1698431365
transform 1 0 161616 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_1437
timestamp 1698431365
transform 1 0 162288 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_1501
timestamp 1698431365
transform 1 0 169456 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_1507
timestamp 1698431365
transform 1 0 170128 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_1571
timestamp 1698431365
transform 1 0 177296 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_1577
timestamp 1698431365
transform 1 0 177968 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_1641
timestamp 1698431365
transform 1 0 185136 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_1647
timestamp 1698431365
transform 1 0 185808 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_1711
timestamp 1698431365
transform 1 0 192976 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_1717
timestamp 1698431365
transform 1 0 193648 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_1781
timestamp 1698431365
transform 1 0 200816 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_1787
timestamp 1698431365
transform 1 0 201488 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_1851
timestamp 1698431365
transform 1 0 208656 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_46_1857
timestamp 1698431365
transform 1 0 209328 0 1 39200
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_1921
timestamp 1698431365
transform 1 0 216496 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_1927
timestamp 1698431365
transform 1 0 217168 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_1935
timestamp 1698431365
transform 1 0 218064 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_1937
timestamp 1698431365
transform 1 0 218288 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_2
timestamp 1698431365
transform 1 0 1568 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_66
timestamp 1698431365
transform 1 0 8736 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_72
timestamp 1698431365
transform 1 0 9408 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_136
timestamp 1698431365
transform 1 0 16576 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_142
timestamp 1698431365
transform 1 0 17248 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_206
timestamp 1698431365
transform 1 0 24416 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_212
timestamp 1698431365
transform 1 0 25088 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_276
timestamp 1698431365
transform 1 0 32256 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_282
timestamp 1698431365
transform 1 0 32928 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_346
timestamp 1698431365
transform 1 0 40096 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_352
timestamp 1698431365
transform 1 0 40768 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_416
timestamp 1698431365
transform 1 0 47936 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_422
timestamp 1698431365
transform 1 0 48608 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_486
timestamp 1698431365
transform 1 0 55776 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_492
timestamp 1698431365
transform 1 0 56448 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_556
timestamp 1698431365
transform 1 0 63616 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_562
timestamp 1698431365
transform 1 0 64288 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_626
timestamp 1698431365
transform 1 0 71456 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_632
timestamp 1698431365
transform 1 0 72128 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_696
timestamp 1698431365
transform 1 0 79296 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_702
timestamp 1698431365
transform 1 0 79968 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_766
timestamp 1698431365
transform 1 0 87136 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_772
timestamp 1698431365
transform 1 0 87808 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_836
timestamp 1698431365
transform 1 0 94976 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_842
timestamp 1698431365
transform 1 0 95648 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_906
timestamp 1698431365
transform 1 0 102816 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_912
timestamp 1698431365
transform 1 0 103488 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_976
timestamp 1698431365
transform 1 0 110656 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_982
timestamp 1698431365
transform 1 0 111328 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_1046
timestamp 1698431365
transform 1 0 118496 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_1052
timestamp 1698431365
transform 1 0 119168 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_1116
timestamp 1698431365
transform 1 0 126336 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_1122
timestamp 1698431365
transform 1 0 127008 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_1186
timestamp 1698431365
transform 1 0 134176 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_1192
timestamp 1698431365
transform 1 0 134848 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_1256
timestamp 1698431365
transform 1 0 142016 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_1262
timestamp 1698431365
transform 1 0 142688 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_1326
timestamp 1698431365
transform 1 0 149856 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_1332
timestamp 1698431365
transform 1 0 150528 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_1396
timestamp 1698431365
transform 1 0 157696 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_1402
timestamp 1698431365
transform 1 0 158368 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_1466
timestamp 1698431365
transform 1 0 165536 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_1472
timestamp 1698431365
transform 1 0 166208 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_1536
timestamp 1698431365
transform 1 0 173376 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_1542
timestamp 1698431365
transform 1 0 174048 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_1606
timestamp 1698431365
transform 1 0 181216 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_1612
timestamp 1698431365
transform 1 0 181888 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_1676
timestamp 1698431365
transform 1 0 189056 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_1682
timestamp 1698431365
transform 1 0 189728 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_1746
timestamp 1698431365
transform 1 0 196896 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_1752
timestamp 1698431365
transform 1 0 197568 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_1816
timestamp 1698431365
transform 1 0 204736 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_47_1822
timestamp 1698431365
transform 1 0 205408 0 -1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_1886
timestamp 1698431365
transform 1 0 212576 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_47_1892
timestamp 1698431365
transform 1 0 213248 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_1924
timestamp 1698431365
transform 1 0 216832 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_1932
timestamp 1698431365
transform 1 0 217728 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_1936
timestamp 1698431365
transform 1 0 218176 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_2
timestamp 1698431365
transform 1 0 1568 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_34
timestamp 1698431365
transform 1 0 5152 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_37
timestamp 1698431365
transform 1 0 5488 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_101
timestamp 1698431365
transform 1 0 12656 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_107
timestamp 1698431365
transform 1 0 13328 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_171
timestamp 1698431365
transform 1 0 20496 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_177
timestamp 1698431365
transform 1 0 21168 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_241
timestamp 1698431365
transform 1 0 28336 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_247
timestamp 1698431365
transform 1 0 29008 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_311
timestamp 1698431365
transform 1 0 36176 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_317
timestamp 1698431365
transform 1 0 36848 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_381
timestamp 1698431365
transform 1 0 44016 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_387
timestamp 1698431365
transform 1 0 44688 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_451
timestamp 1698431365
transform 1 0 51856 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_457
timestamp 1698431365
transform 1 0 52528 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_521
timestamp 1698431365
transform 1 0 59696 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_527
timestamp 1698431365
transform 1 0 60368 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_591
timestamp 1698431365
transform 1 0 67536 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_597
timestamp 1698431365
transform 1 0 68208 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_661
timestamp 1698431365
transform 1 0 75376 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_667
timestamp 1698431365
transform 1 0 76048 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_731
timestamp 1698431365
transform 1 0 83216 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_737
timestamp 1698431365
transform 1 0 83888 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_801
timestamp 1698431365
transform 1 0 91056 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_807
timestamp 1698431365
transform 1 0 91728 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_871
timestamp 1698431365
transform 1 0 98896 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_877
timestamp 1698431365
transform 1 0 99568 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_941
timestamp 1698431365
transform 1 0 106736 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_947
timestamp 1698431365
transform 1 0 107408 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_1011
timestamp 1698431365
transform 1 0 114576 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_1017
timestamp 1698431365
transform 1 0 115248 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_1081
timestamp 1698431365
transform 1 0 122416 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_1087
timestamp 1698431365
transform 1 0 123088 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_1151
timestamp 1698431365
transform 1 0 130256 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_1157
timestamp 1698431365
transform 1 0 130928 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_1221
timestamp 1698431365
transform 1 0 138096 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_1227
timestamp 1698431365
transform 1 0 138768 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_1291
timestamp 1698431365
transform 1 0 145936 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_1297
timestamp 1698431365
transform 1 0 146608 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_1361
timestamp 1698431365
transform 1 0 153776 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_1367
timestamp 1698431365
transform 1 0 154448 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_1431
timestamp 1698431365
transform 1 0 161616 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_1437
timestamp 1698431365
transform 1 0 162288 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_1501
timestamp 1698431365
transform 1 0 169456 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_1507
timestamp 1698431365
transform 1 0 170128 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_1571
timestamp 1698431365
transform 1 0 177296 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_1577
timestamp 1698431365
transform 1 0 177968 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_1641
timestamp 1698431365
transform 1 0 185136 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_1647
timestamp 1698431365
transform 1 0 185808 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_1711
timestamp 1698431365
transform 1 0 192976 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_1717
timestamp 1698431365
transform 1 0 193648 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_1781
timestamp 1698431365
transform 1 0 200816 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_1787
timestamp 1698431365
transform 1 0 201488 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_1851
timestamp 1698431365
transform 1 0 208656 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_1857
timestamp 1698431365
transform 1 0 209328 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_1921
timestamp 1698431365
transform 1 0 216496 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_1927
timestamp 1698431365
transform 1 0 217168 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_1935
timestamp 1698431365
transform 1 0 218064 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_1937
timestamp 1698431365
transform 1 0 218288 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_2
timestamp 1698431365
transform 1 0 1568 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_66
timestamp 1698431365
transform 1 0 8736 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_72
timestamp 1698431365
transform 1 0 9408 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_136
timestamp 1698431365
transform 1 0 16576 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_142
timestamp 1698431365
transform 1 0 17248 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_206
timestamp 1698431365
transform 1 0 24416 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_212
timestamp 1698431365
transform 1 0 25088 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_276
timestamp 1698431365
transform 1 0 32256 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_282
timestamp 1698431365
transform 1 0 32928 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_346
timestamp 1698431365
transform 1 0 40096 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_352
timestamp 1698431365
transform 1 0 40768 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_416
timestamp 1698431365
transform 1 0 47936 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_422
timestamp 1698431365
transform 1 0 48608 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_486
timestamp 1698431365
transform 1 0 55776 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_492
timestamp 1698431365
transform 1 0 56448 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_556
timestamp 1698431365
transform 1 0 63616 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_562
timestamp 1698431365
transform 1 0 64288 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_626
timestamp 1698431365
transform 1 0 71456 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_632
timestamp 1698431365
transform 1 0 72128 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_696
timestamp 1698431365
transform 1 0 79296 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_702
timestamp 1698431365
transform 1 0 79968 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_766
timestamp 1698431365
transform 1 0 87136 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_772
timestamp 1698431365
transform 1 0 87808 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_836
timestamp 1698431365
transform 1 0 94976 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_842
timestamp 1698431365
transform 1 0 95648 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_906
timestamp 1698431365
transform 1 0 102816 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_912
timestamp 1698431365
transform 1 0 103488 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_976
timestamp 1698431365
transform 1 0 110656 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_982
timestamp 1698431365
transform 1 0 111328 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_1046
timestamp 1698431365
transform 1 0 118496 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_1052
timestamp 1698431365
transform 1 0 119168 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_1116
timestamp 1698431365
transform 1 0 126336 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_1122
timestamp 1698431365
transform 1 0 127008 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_1186
timestamp 1698431365
transform 1 0 134176 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_1192
timestamp 1698431365
transform 1 0 134848 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_1256
timestamp 1698431365
transform 1 0 142016 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_1262
timestamp 1698431365
transform 1 0 142688 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_1326
timestamp 1698431365
transform 1 0 149856 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_1332
timestamp 1698431365
transform 1 0 150528 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_1396
timestamp 1698431365
transform 1 0 157696 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_1402
timestamp 1698431365
transform 1 0 158368 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_1466
timestamp 1698431365
transform 1 0 165536 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_1472
timestamp 1698431365
transform 1 0 166208 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_1536
timestamp 1698431365
transform 1 0 173376 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_1542
timestamp 1698431365
transform 1 0 174048 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_1606
timestamp 1698431365
transform 1 0 181216 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_1612
timestamp 1698431365
transform 1 0 181888 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_1676
timestamp 1698431365
transform 1 0 189056 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_1682
timestamp 1698431365
transform 1 0 189728 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_1746
timestamp 1698431365
transform 1 0 196896 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_1752
timestamp 1698431365
transform 1 0 197568 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_1816
timestamp 1698431365
transform 1 0 204736 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_49_1822
timestamp 1698431365
transform 1 0 205408 0 -1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_1886
timestamp 1698431365
transform 1 0 212576 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_1892
timestamp 1698431365
transform 1 0 213248 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_1924
timestamp 1698431365
transform 1 0 216832 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_1932
timestamp 1698431365
transform 1 0 217728 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_1936
timestamp 1698431365
transform 1 0 218176 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_2
timestamp 1698431365
transform 1 0 1568 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_34
timestamp 1698431365
transform 1 0 5152 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_37
timestamp 1698431365
transform 1 0 5488 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_101
timestamp 1698431365
transform 1 0 12656 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_107
timestamp 1698431365
transform 1 0 13328 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_171
timestamp 1698431365
transform 1 0 20496 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_177
timestamp 1698431365
transform 1 0 21168 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_241
timestamp 1698431365
transform 1 0 28336 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_247
timestamp 1698431365
transform 1 0 29008 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_311
timestamp 1698431365
transform 1 0 36176 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_317
timestamp 1698431365
transform 1 0 36848 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_381
timestamp 1698431365
transform 1 0 44016 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_387
timestamp 1698431365
transform 1 0 44688 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_451
timestamp 1698431365
transform 1 0 51856 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_457
timestamp 1698431365
transform 1 0 52528 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_521
timestamp 1698431365
transform 1 0 59696 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_527
timestamp 1698431365
transform 1 0 60368 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_591
timestamp 1698431365
transform 1 0 67536 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_597
timestamp 1698431365
transform 1 0 68208 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_661
timestamp 1698431365
transform 1 0 75376 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_667
timestamp 1698431365
transform 1 0 76048 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_731
timestamp 1698431365
transform 1 0 83216 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_737
timestamp 1698431365
transform 1 0 83888 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_801
timestamp 1698431365
transform 1 0 91056 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_807
timestamp 1698431365
transform 1 0 91728 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_871
timestamp 1698431365
transform 1 0 98896 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_877
timestamp 1698431365
transform 1 0 99568 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_941
timestamp 1698431365
transform 1 0 106736 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_947
timestamp 1698431365
transform 1 0 107408 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_1011
timestamp 1698431365
transform 1 0 114576 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_1017
timestamp 1698431365
transform 1 0 115248 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_1081
timestamp 1698431365
transform 1 0 122416 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_1087
timestamp 1698431365
transform 1 0 123088 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_1151
timestamp 1698431365
transform 1 0 130256 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_1157
timestamp 1698431365
transform 1 0 130928 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_1189
timestamp 1698431365
transform 1 0 134512 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_1205
timestamp 1698431365
transform 1 0 136304 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_1213
timestamp 1698431365
transform 1 0 137200 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_1215
timestamp 1698431365
transform 1 0 137424 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_1224
timestamp 1698431365
transform 1 0 138432 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_1227
timestamp 1698431365
transform 1 0 138768 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_1291
timestamp 1698431365
transform 1 0 145936 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_1297
timestamp 1698431365
transform 1 0 146608 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_1361
timestamp 1698431365
transform 1 0 153776 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_1367
timestamp 1698431365
transform 1 0 154448 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_1431
timestamp 1698431365
transform 1 0 161616 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_1437
timestamp 1698431365
transform 1 0 162288 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_1501
timestamp 1698431365
transform 1 0 169456 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_1507
timestamp 1698431365
transform 1 0 170128 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_1571
timestamp 1698431365
transform 1 0 177296 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_1577
timestamp 1698431365
transform 1 0 177968 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_1641
timestamp 1698431365
transform 1 0 185136 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_1647
timestamp 1698431365
transform 1 0 185808 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_1711
timestamp 1698431365
transform 1 0 192976 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_1717
timestamp 1698431365
transform 1 0 193648 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_1781
timestamp 1698431365
transform 1 0 200816 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_1787
timestamp 1698431365
transform 1 0 201488 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_1851
timestamp 1698431365
transform 1 0 208656 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_50_1857
timestamp 1698431365
transform 1 0 209328 0 1 42336
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_1921
timestamp 1698431365
transform 1 0 216496 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_1927
timestamp 1698431365
transform 1 0 217168 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_1935
timestamp 1698431365
transform 1 0 218064 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_1937
timestamp 1698431365
transform 1 0 218288 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_2
timestamp 1698431365
transform 1 0 1568 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_66
timestamp 1698431365
transform 1 0 8736 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_72
timestamp 1698431365
transform 1 0 9408 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_136
timestamp 1698431365
transform 1 0 16576 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_142
timestamp 1698431365
transform 1 0 17248 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_206
timestamp 1698431365
transform 1 0 24416 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_212
timestamp 1698431365
transform 1 0 25088 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_276
timestamp 1698431365
transform 1 0 32256 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_282
timestamp 1698431365
transform 1 0 32928 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_346
timestamp 1698431365
transform 1 0 40096 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_352
timestamp 1698431365
transform 1 0 40768 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_416
timestamp 1698431365
transform 1 0 47936 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_422
timestamp 1698431365
transform 1 0 48608 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_486
timestamp 1698431365
transform 1 0 55776 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_492
timestamp 1698431365
transform 1 0 56448 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_556
timestamp 1698431365
transform 1 0 63616 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_562
timestamp 1698431365
transform 1 0 64288 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_626
timestamp 1698431365
transform 1 0 71456 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_632
timestamp 1698431365
transform 1 0 72128 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_696
timestamp 1698431365
transform 1 0 79296 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_702
timestamp 1698431365
transform 1 0 79968 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_766
timestamp 1698431365
transform 1 0 87136 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_772
timestamp 1698431365
transform 1 0 87808 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_836
timestamp 1698431365
transform 1 0 94976 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_842
timestamp 1698431365
transform 1 0 95648 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_906
timestamp 1698431365
transform 1 0 102816 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_912
timestamp 1698431365
transform 1 0 103488 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_976
timestamp 1698431365
transform 1 0 110656 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_982
timestamp 1698431365
transform 1 0 111328 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_1046
timestamp 1698431365
transform 1 0 118496 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_1052
timestamp 1698431365
transform 1 0 119168 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_1116
timestamp 1698431365
transform 1 0 126336 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_1122
timestamp 1698431365
transform 1 0 127008 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_1186
timestamp 1698431365
transform 1 0 134176 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_1192
timestamp 1698431365
transform 1 0 134848 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_1196
timestamp 1698431365
transform 1 0 135296 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_1198
timestamp 1698431365
transform 1 0 135520 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_1206
timestamp 1698431365
transform 1 0 136416 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_1210
timestamp 1698431365
transform 1 0 136864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_1212
timestamp 1698431365
transform 1 0 137088 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_1244
timestamp 1698431365
transform 1 0 140672 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_1262
timestamp 1698431365
transform 1 0 142688 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_1326
timestamp 1698431365
transform 1 0 149856 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_1332
timestamp 1698431365
transform 1 0 150528 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_1396
timestamp 1698431365
transform 1 0 157696 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_1402
timestamp 1698431365
transform 1 0 158368 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_1466
timestamp 1698431365
transform 1 0 165536 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_1472
timestamp 1698431365
transform 1 0 166208 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_1536
timestamp 1698431365
transform 1 0 173376 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_1542
timestamp 1698431365
transform 1 0 174048 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_1606
timestamp 1698431365
transform 1 0 181216 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_1612
timestamp 1698431365
transform 1 0 181888 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_1676
timestamp 1698431365
transform 1 0 189056 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_1682
timestamp 1698431365
transform 1 0 189728 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_1746
timestamp 1698431365
transform 1 0 196896 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_1752
timestamp 1698431365
transform 1 0 197568 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_1816
timestamp 1698431365
transform 1 0 204736 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_1822
timestamp 1698431365
transform 1 0 205408 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_1886
timestamp 1698431365
transform 1 0 212576 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_51_1892
timestamp 1698431365
transform 1 0 213248 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_1924
timestamp 1698431365
transform 1 0 216832 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_1932
timestamp 1698431365
transform 1 0 217728 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_1936
timestamp 1698431365
transform 1 0 218176 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_2
timestamp 1698431365
transform 1 0 1568 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_34
timestamp 1698431365
transform 1 0 5152 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_37
timestamp 1698431365
transform 1 0 5488 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_101
timestamp 1698431365
transform 1 0 12656 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_107
timestamp 1698431365
transform 1 0 13328 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_171
timestamp 1698431365
transform 1 0 20496 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_177
timestamp 1698431365
transform 1 0 21168 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_241
timestamp 1698431365
transform 1 0 28336 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_247
timestamp 1698431365
transform 1 0 29008 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_311
timestamp 1698431365
transform 1 0 36176 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_317
timestamp 1698431365
transform 1 0 36848 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_381
timestamp 1698431365
transform 1 0 44016 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_387
timestamp 1698431365
transform 1 0 44688 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_451
timestamp 1698431365
transform 1 0 51856 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_457
timestamp 1698431365
transform 1 0 52528 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_521
timestamp 1698431365
transform 1 0 59696 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_527
timestamp 1698431365
transform 1 0 60368 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_591
timestamp 1698431365
transform 1 0 67536 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_597
timestamp 1698431365
transform 1 0 68208 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_661
timestamp 1698431365
transform 1 0 75376 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_667
timestamp 1698431365
transform 1 0 76048 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_731
timestamp 1698431365
transform 1 0 83216 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_737
timestamp 1698431365
transform 1 0 83888 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_801
timestamp 1698431365
transform 1 0 91056 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_807
timestamp 1698431365
transform 1 0 91728 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_871
timestamp 1698431365
transform 1 0 98896 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_877
timestamp 1698431365
transform 1 0 99568 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_941
timestamp 1698431365
transform 1 0 106736 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_947
timestamp 1698431365
transform 1 0 107408 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_1011
timestamp 1698431365
transform 1 0 114576 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_1017
timestamp 1698431365
transform 1 0 115248 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_1081
timestamp 1698431365
transform 1 0 122416 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_1087
timestamp 1698431365
transform 1 0 123088 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_1151
timestamp 1698431365
transform 1 0 130256 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_1157
timestamp 1698431365
transform 1 0 130928 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_1161
timestamp 1698431365
transform 1 0 131376 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_1163
timestamp 1698431365
transform 1 0 131600 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_1222
timestamp 1698431365
transform 1 0 138208 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_1224
timestamp 1698431365
transform 1 0 138432 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_1256
timestamp 1698431365
transform 1 0 142016 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_1288
timestamp 1698431365
transform 1 0 145600 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_1292
timestamp 1698431365
transform 1 0 146048 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_1294
timestamp 1698431365
transform 1 0 146272 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_1297
timestamp 1698431365
transform 1 0 146608 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_1361
timestamp 1698431365
transform 1 0 153776 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_1367
timestamp 1698431365
transform 1 0 154448 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_1431
timestamp 1698431365
transform 1 0 161616 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_1437
timestamp 1698431365
transform 1 0 162288 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_1501
timestamp 1698431365
transform 1 0 169456 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_1507
timestamp 1698431365
transform 1 0 170128 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_1571
timestamp 1698431365
transform 1 0 177296 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_1577
timestamp 1698431365
transform 1 0 177968 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_1641
timestamp 1698431365
transform 1 0 185136 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_1647
timestamp 1698431365
transform 1 0 185808 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_1711
timestamp 1698431365
transform 1 0 192976 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_1717
timestamp 1698431365
transform 1 0 193648 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_1781
timestamp 1698431365
transform 1 0 200816 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_1787
timestamp 1698431365
transform 1 0 201488 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_1851
timestamp 1698431365
transform 1 0 208656 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_52_1857
timestamp 1698431365
transform 1 0 209328 0 1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_1921
timestamp 1698431365
transform 1 0 216496 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_1927
timestamp 1698431365
transform 1 0 217168 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_1935
timestamp 1698431365
transform 1 0 218064 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_1937
timestamp 1698431365
transform 1 0 218288 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_2
timestamp 1698431365
transform 1 0 1568 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_66
timestamp 1698431365
transform 1 0 8736 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_72
timestamp 1698431365
transform 1 0 9408 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_136
timestamp 1698431365
transform 1 0 16576 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_142
timestamp 1698431365
transform 1 0 17248 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_206
timestamp 1698431365
transform 1 0 24416 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_212
timestamp 1698431365
transform 1 0 25088 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_276
timestamp 1698431365
transform 1 0 32256 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_282
timestamp 1698431365
transform 1 0 32928 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_346
timestamp 1698431365
transform 1 0 40096 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_352
timestamp 1698431365
transform 1 0 40768 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_416
timestamp 1698431365
transform 1 0 47936 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_422
timestamp 1698431365
transform 1 0 48608 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_486
timestamp 1698431365
transform 1 0 55776 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_492
timestamp 1698431365
transform 1 0 56448 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_556
timestamp 1698431365
transform 1 0 63616 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_562
timestamp 1698431365
transform 1 0 64288 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_626
timestamp 1698431365
transform 1 0 71456 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_632
timestamp 1698431365
transform 1 0 72128 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_648
timestamp 1698431365
transform 1 0 73920 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_656
timestamp 1698431365
transform 1 0 74816 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_660
timestamp 1698431365
transform 1 0 75264 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_662
timestamp 1698431365
transform 1 0 75488 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_689
timestamp 1698431365
transform 1 0 78512 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_693
timestamp 1698431365
transform 1 0 78960 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_697
timestamp 1698431365
transform 1 0 79408 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_699
timestamp 1698431365
transform 1 0 79632 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_702
timestamp 1698431365
transform 1 0 79968 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_766
timestamp 1698431365
transform 1 0 87136 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_772
timestamp 1698431365
transform 1 0 87808 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_836
timestamp 1698431365
transform 1 0 94976 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_842
timestamp 1698431365
transform 1 0 95648 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_906
timestamp 1698431365
transform 1 0 102816 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_912
timestamp 1698431365
transform 1 0 103488 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_976
timestamp 1698431365
transform 1 0 110656 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_982
timestamp 1698431365
transform 1 0 111328 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_1046
timestamp 1698431365
transform 1 0 118496 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_1052
timestamp 1698431365
transform 1 0 119168 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_1116
timestamp 1698431365
transform 1 0 126336 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_1122
timestamp 1698431365
transform 1 0 127008 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_1186
timestamp 1698431365
transform 1 0 134176 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_1192
timestamp 1698431365
transform 1 0 134848 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_1196
timestamp 1698431365
transform 1 0 135296 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_1212
timestamp 1698431365
transform 1 0 137088 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_1220
timestamp 1698431365
transform 1 0 137984 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_1223
timestamp 1698431365
transform 1 0 138320 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_1227
timestamp 1698431365
transform 1 0 138768 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_1254
timestamp 1698431365
transform 1 0 141792 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_1258
timestamp 1698431365
transform 1 0 142240 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_1262
timestamp 1698431365
transform 1 0 142688 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_1326
timestamp 1698431365
transform 1 0 149856 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_1332
timestamp 1698431365
transform 1 0 150528 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_1340
timestamp 1698431365
transform 1 0 151424 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_1344
timestamp 1698431365
transform 1 0 151872 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_1373
timestamp 1698431365
transform 1 0 155120 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_1389
timestamp 1698431365
transform 1 0 156912 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_1397
timestamp 1698431365
transform 1 0 157808 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_1399
timestamp 1698431365
transform 1 0 158032 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_1402
timestamp 1698431365
transform 1 0 158368 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_1466
timestamp 1698431365
transform 1 0 165536 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_1472
timestamp 1698431365
transform 1 0 166208 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_1536
timestamp 1698431365
transform 1 0 173376 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_1542
timestamp 1698431365
transform 1 0 174048 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_1606
timestamp 1698431365
transform 1 0 181216 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_1612
timestamp 1698431365
transform 1 0 181888 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_1676
timestamp 1698431365
transform 1 0 189056 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_1682
timestamp 1698431365
transform 1 0 189728 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_1746
timestamp 1698431365
transform 1 0 196896 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_1752
timestamp 1698431365
transform 1 0 197568 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_1816
timestamp 1698431365
transform 1 0 204736 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_1822
timestamp 1698431365
transform 1 0 205408 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_1886
timestamp 1698431365
transform 1 0 212576 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_53_1892
timestamp 1698431365
transform 1 0 213248 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_1924
timestamp 1698431365
transform 1 0 216832 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_1932
timestamp 1698431365
transform 1 0 217728 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_1936
timestamp 1698431365
transform 1 0 218176 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_2
timestamp 1698431365
transform 1 0 1568 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_36
timestamp 1698431365
transform 1 0 5376 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_44
timestamp 1698431365
transform 1 0 6272 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_48
timestamp 1698431365
transform 1 0 6720 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_57
timestamp 1698431365
transform 1 0 7728 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_65
timestamp 1698431365
transform 1 0 8624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_67
timestamp 1698431365
transform 1 0 8848 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_70
timestamp 1698431365
transform 1 0 9184 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_78
timestamp 1698431365
transform 1 0 10080 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_82
timestamp 1698431365
transform 1 0 10528 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_84
timestamp 1698431365
transform 1 0 10752 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_101
timestamp 1698431365
transform 1 0 12656 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_104
timestamp 1698431365
transform 1 0 12992 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_120
timestamp 1698431365
transform 1 0 14784 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_131
timestamp 1698431365
transform 1 0 16016 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_135
timestamp 1698431365
transform 1 0 16464 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_138
timestamp 1698431365
transform 1 0 16800 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_154
timestamp 1698431365
transform 1 0 18592 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_156
timestamp 1698431365
transform 1 0 18816 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_167
timestamp 1698431365
transform 1 0 20048 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_169
timestamp 1698431365
transform 1 0 20272 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_172
timestamp 1698431365
transform 1 0 20608 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_188
timestamp 1698431365
transform 1 0 22400 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_192
timestamp 1698431365
transform 1 0 22848 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_203
timestamp 1698431365
transform 1 0 24080 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_206
timestamp 1698431365
transform 1 0 24416 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_222
timestamp 1698431365
transform 1 0 26208 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_230
timestamp 1698431365
transform 1 0 27104 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_234
timestamp 1698431365
transform 1 0 27552 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_248
timestamp 1698431365
transform 1 0 29120 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_264
timestamp 1698431365
transform 1 0 30912 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_268
timestamp 1698431365
transform 1 0 31360 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_282
timestamp 1698431365
transform 1 0 32928 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_298
timestamp 1698431365
transform 1 0 34720 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_302
timestamp 1698431365
transform 1 0 35168 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_316
timestamp 1698431365
transform 1 0 36736 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_332
timestamp 1698431365
transform 1 0 38528 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_336
timestamp 1698431365
transform 1 0 38976 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_350
timestamp 1698431365
transform 1 0 40544 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_366
timestamp 1698431365
transform 1 0 42336 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_370
timestamp 1698431365
transform 1 0 42784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_384
timestamp 1698431365
transform 1 0 44352 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_400
timestamp 1698431365
transform 1 0 46144 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_410
timestamp 1698431365
transform 1 0 47264 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_437
timestamp 1698431365
transform 1 0 50288 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_441
timestamp 1698431365
transform 1 0 50736 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_444
timestamp 1698431365
transform 1 0 51072 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_446
timestamp 1698431365
transform 1 0 51296 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_473
timestamp 1698431365
transform 1 0 54320 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_475
timestamp 1698431365
transform 1 0 54544 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_478
timestamp 1698431365
transform 1 0 54880 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_482
timestamp 1698431365
transform 1 0 55328 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_509
timestamp 1698431365
transform 1 0 58352 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_512
timestamp 1698431365
transform 1 0 58688 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_516
timestamp 1698431365
transform 1 0 59136 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_546
timestamp 1698431365
transform 1 0 62496 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_550
timestamp 1698431365
transform 1 0 62944 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_580
timestamp 1698431365
transform 1 0 66304 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_584
timestamp 1698431365
transform 1 0 66752 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_614
timestamp 1698431365
transform 1 0 70112 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_618
timestamp 1698431365
transform 1 0 70560 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_648
timestamp 1698431365
transform 1 0 73920 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_652
timestamp 1698431365
transform 1 0 74368 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_668
timestamp 1698431365
transform 1 0 76160 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_676
timestamp 1698431365
transform 1 0 77056 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_682
timestamp 1698431365
transform 1 0 77728 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_690
timestamp 1698431365
transform 1 0 78624 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_694
timestamp 1698431365
transform 1 0 79072 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_696
timestamp 1698431365
transform 1 0 79296 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_705
timestamp 1698431365
transform 1 0 80304 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_713
timestamp 1698431365
transform 1 0 81200 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_716
timestamp 1698431365
transform 1 0 81536 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_732
timestamp 1698431365
transform 1 0 83328 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_741
timestamp 1698431365
transform 1 0 84336 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_745
timestamp 1698431365
transform 1 0 84784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_747
timestamp 1698431365
transform 1 0 85008 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_750
timestamp 1698431365
transform 1 0 85344 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_766
timestamp 1698431365
transform 1 0 87136 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_768
timestamp 1698431365
transform 1 0 87360 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_777
timestamp 1698431365
transform 1 0 88368 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_781
timestamp 1698431365
transform 1 0 88816 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_784
timestamp 1698431365
transform 1 0 89152 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_800
timestamp 1698431365
transform 1 0 90944 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_804
timestamp 1698431365
transform 1 0 91392 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_813
timestamp 1698431365
transform 1 0 92400 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_815
timestamp 1698431365
transform 1 0 92624 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_818
timestamp 1698431365
transform 1 0 92960 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_834
timestamp 1698431365
transform 1 0 94752 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_838
timestamp 1698431365
transform 1 0 95200 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_840
timestamp 1698431365
transform 1 0 95424 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_849
timestamp 1698431365
transform 1 0 96432 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_852
timestamp 1698431365
transform 1 0 96768 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_868
timestamp 1698431365
transform 1 0 98560 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_876
timestamp 1698431365
transform 1 0 99456 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_880
timestamp 1698431365
transform 1 0 99904 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_892
timestamp 1698431365
transform 1 0 101248 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_908
timestamp 1698431365
transform 1 0 103040 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_926
timestamp 1698431365
transform 1 0 105056 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_942
timestamp 1698431365
transform 1 0 106848 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_960
timestamp 1698431365
transform 1 0 108864 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_976
timestamp 1698431365
transform 1 0 110656 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_994
timestamp 1698431365
transform 1 0 112672 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_1010
timestamp 1698431365
transform 1 0 114464 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_1022
timestamp 1698431365
transform 1 0 115808 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_1029
timestamp 1698431365
transform 1 0 116592 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_1045
timestamp 1698431365
transform 1 0 118384 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_1049
timestamp 1698431365
transform 1 0 118832 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_1051
timestamp 1698431365
transform 1 0 119056 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_1056
timestamp 1698431365
transform 1 0 119616 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_1058
timestamp 1698431365
transform 1 0 119840 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_1065
timestamp 1698431365
transform 1 0 120624 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_1081
timestamp 1698431365
transform 1 0 122416 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_1085
timestamp 1698431365
transform 1 0 122864 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_1087
timestamp 1698431365
transform 1 0 123088 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_1090
timestamp 1698431365
transform 1 0 123424 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_1092
timestamp 1698431365
transform 1 0 123648 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_1101
timestamp 1698431365
transform 1 0 124656 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_1117
timestamp 1698431365
transform 1 0 126448 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_1121
timestamp 1698431365
transform 1 0 126896 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_1124
timestamp 1698431365
transform 1 0 127232 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_1128
timestamp 1698431365
transform 1 0 127680 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_1137
timestamp 1698431365
transform 1 0 128688 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_1153
timestamp 1698431365
transform 1 0 130480 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_1155
timestamp 1698431365
transform 1 0 130704 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_1158
timestamp 1698431365
transform 1 0 131040 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_1162
timestamp 1698431365
transform 1 0 131488 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_1164
timestamp 1698431365
transform 1 0 131712 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_1173
timestamp 1698431365
transform 1 0 132720 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_1189
timestamp 1698431365
transform 1 0 134512 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_1192
timestamp 1698431365
transform 1 0 134848 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_1200
timestamp 1698431365
transform 1 0 135744 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_1209
timestamp 1698431365
transform 1 0 136752 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_1217
timestamp 1698431365
transform 1 0 137648 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_1221
timestamp 1698431365
transform 1 0 138096 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_1223
timestamp 1698431365
transform 1 0 138320 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_1226
timestamp 1698431365
transform 1 0 138656 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_1234
timestamp 1698431365
transform 1 0 139552 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_1236
timestamp 1698431365
transform 1 0 139776 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_1245
timestamp 1698431365
transform 1 0 140784 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_1253
timestamp 1698431365
transform 1 0 141680 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_1257
timestamp 1698431365
transform 1 0 142128 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_1260
timestamp 1698431365
transform 1 0 142464 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_1268
timestamp 1698431365
transform 1 0 143360 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_1272
timestamp 1698431365
transform 1 0 143808 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_1281
timestamp 1698431365
transform 1 0 144816 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_1289
timestamp 1698431365
transform 1 0 145712 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_1291
timestamp 1698431365
transform 1 0 145936 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_1294
timestamp 1698431365
transform 1 0 146272 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_1354
timestamp 1698431365
transform 1 0 152992 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_1358
timestamp 1698431365
transform 1 0 153440 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_1362
timestamp 1698431365
transform 1 0 153888 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_1378
timestamp 1698431365
transform 1 0 155680 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_1380
timestamp 1698431365
transform 1 0 155904 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_1389
timestamp 1698431365
transform 1 0 156912 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_1393
timestamp 1698431365
transform 1 0 157360 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_1396
timestamp 1698431365
transform 1 0 157696 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_1412
timestamp 1698431365
transform 1 0 159488 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_1416
timestamp 1698431365
transform 1 0 159936 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_1425
timestamp 1698431365
transform 1 0 160944 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_1427
timestamp 1698431365
transform 1 0 161168 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_1430
timestamp 1698431365
transform 1 0 161504 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_1446
timestamp 1698431365
transform 1 0 163296 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_1450
timestamp 1698431365
transform 1 0 163744 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_1452
timestamp 1698431365
transform 1 0 163968 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_1461
timestamp 1698431365
transform 1 0 164976 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_1464
timestamp 1698431365
transform 1 0 165312 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_1480
timestamp 1698431365
transform 1 0 167104 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_1488
timestamp 1698431365
transform 1 0 168000 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_1492
timestamp 1698431365
transform 1 0 168448 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_1504
timestamp 1698431365
transform 1 0 169792 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_1520
timestamp 1698431365
transform 1 0 171584 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_1538
timestamp 1698431365
transform 1 0 173600 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_1554
timestamp 1698431365
transform 1 0 175392 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_1572
timestamp 1698431365
transform 1 0 177408 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_1588
timestamp 1698431365
transform 1 0 179200 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_1606
timestamp 1698431365
transform 1 0 181216 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_1622
timestamp 1698431365
transform 1 0 183008 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_1634
timestamp 1698431365
transform 1 0 184352 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_1641
timestamp 1698431365
transform 1 0 185136 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_1657
timestamp 1698431365
transform 1 0 186928 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_1661
timestamp 1698431365
transform 1 0 187376 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_1663
timestamp 1698431365
transform 1 0 187600 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_1668
timestamp 1698431365
transform 1 0 188160 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_1670
timestamp 1698431365
transform 1 0 188384 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_1679
timestamp 1698431365
transform 1 0 189392 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_1695
timestamp 1698431365
transform 1 0 191184 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_1699
timestamp 1698431365
transform 1 0 191632 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_1702
timestamp 1698431365
transform 1 0 191968 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_1704
timestamp 1698431365
transform 1 0 192192 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_1715
timestamp 1698431365
transform 1 0 193424 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_1731
timestamp 1698431365
transform 1 0 195216 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_1733
timestamp 1698431365
transform 1 0 195440 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_1736
timestamp 1698431365
transform 1 0 195776 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_1740
timestamp 1698431365
transform 1 0 196224 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_1751
timestamp 1698431365
transform 1 0 197456 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_1767
timestamp 1698431365
transform 1 0 199248 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_1770
timestamp 1698431365
transform 1 0 199584 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_1774
timestamp 1698431365
transform 1 0 200032 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_1776
timestamp 1698431365
transform 1 0 200256 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_1787
timestamp 1698431365
transform 1 0 201488 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_1795
timestamp 1698431365
transform 1 0 202384 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_1799
timestamp 1698431365
transform 1 0 202832 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_1801
timestamp 1698431365
transform 1 0 203056 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_1804
timestamp 1698431365
transform 1 0 203392 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_1812
timestamp 1698431365
transform 1 0 204288 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_1823
timestamp 1698431365
transform 1 0 205520 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_1831
timestamp 1698431365
transform 1 0 206416 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_1835
timestamp 1698431365
transform 1 0 206864 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_1838
timestamp 1698431365
transform 1 0 207200 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_1846
timestamp 1698431365
transform 1 0 208096 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_1848
timestamp 1698431365
transform 1 0 208320 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_1859
timestamp 1698431365
transform 1 0 209552 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_1867
timestamp 1698431365
transform 1 0 210448 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_1869
timestamp 1698431365
transform 1 0 210672 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_1872
timestamp 1698431365
transform 1 0 211008 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_1880
timestamp 1698431365
transform 1 0 211904 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_1884
timestamp 1698431365
transform 1 0 212352 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_1901
timestamp 1698431365
transform 1 0 214256 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_1903
timestamp 1698431365
transform 1 0 214480 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_1906
timestamp 1698431365
transform 1 0 214816 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_1914
timestamp 1698431365
transform 1 0 215712 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_1918
timestamp 1698431365
transform 1 0 216160 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_1920
timestamp 1698431365
transform 1 0 216384 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_1937
timestamp 1698431365
transform 1 0 218288 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input1
timestamp 1698431365
transform 1 0 89712 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input2
timestamp 1698431365
transform 1 0 92960 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input3
timestamp 1698431365
transform 1 0 95088 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698431365
transform 1 0 97776 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform 1 0 100576 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform 1 0 103152 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698431365
transform 1 0 105840 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1698431365
transform 1 0 108528 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input9
timestamp 1698431365
transform 1 0 112000 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1698431365
transform 1 0 113904 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1698431365
transform 1 0 116592 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1698431365
transform 1 0 119616 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1698431365
transform 1 0 121968 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input14
timestamp 1698431365
transform 1 0 124656 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input15
timestamp 1698431365
transform 1 0 127344 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input16
timestamp 1698431365
transform 1 0 130032 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input17
timestamp 1698431365
transform 1 0 132720 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input18
timestamp 1698431365
transform 1 0 135408 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input19
timestamp 1698431365
transform 1 0 138656 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input20
timestamp 1698431365
transform 1 0 140784 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input21
timestamp 1698431365
transform 1 0 143472 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input22
timestamp 1698431365
transform 1 0 146272 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input23
timestamp 1698431365
transform 1 0 148848 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input24
timestamp 1698431365
transform -1 0 153552 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input25
timestamp 1698431365
transform 1 0 154784 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input26
timestamp 1698431365
transform -1 0 158368 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input27
timestamp 1698431365
transform -1 0 160272 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input28
timestamp 1698431365
transform -1 0 163856 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input29
timestamp 1698431365
transform -1 0 165984 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input30
timestamp 1698431365
transform -1 0 168336 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input31
timestamp 1698431365
transform -1 0 171024 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input32
timestamp 1698431365
transform -1 0 173712 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input33
timestamp 1698431365
transform -1 0 176400 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input34
timestamp 1698431365
transform -1 0 179088 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input35
timestamp 1698431365
transform -1 0 181776 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input36
timestamp 1698431365
transform -1 0 185024 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input37
timestamp 1698431365
transform -1 0 187152 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input38
timestamp 1698431365
transform -1 0 189840 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input39
timestamp 1698431365
transform -1 0 192640 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input40
timestamp 1698431365
transform -1 0 195216 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input41
timestamp 1698431365
transform 1 0 197232 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input42
timestamp 1698431365
transform 1 0 199920 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input43
timestamp 1698431365
transform 1 0 203392 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input44
timestamp 1698431365
transform 1 0 205296 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input45
timestamp 1698431365
transform 1 0 207984 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input46
timestamp 1698431365
transform 1 0 211008 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input47
timestamp 1698431365
transform 1 0 213360 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input48
timestamp 1698431365
transform 1 0 216048 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input49
timestamp 1698431365
transform 1 0 156240 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input50
timestamp 1698431365
transform -1 0 160944 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input51
timestamp 1698431365
transform -1 0 164976 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input52
timestamp 1698431365
transform -1 0 169792 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input53
timestamp 1698431365
transform -1 0 173600 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input54
timestamp 1698431365
transform -1 0 177408 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input55
timestamp 1698431365
transform -1 0 181216 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input56
timestamp 1698431365
transform -1 0 185136 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input57
timestamp 1698431365
transform 1 0 188496 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input58
timestamp 1698431365
transform 1 0 192528 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input59
timestamp 1698431365
transform 1 0 196560 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input60
timestamp 1698431365
transform 1 0 200592 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input61
timestamp 1698431365
transform 1 0 204624 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  input62
timestamp 1698431365
transform 1 0 208656 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  input63
timestamp 1698431365
transform 1 0 212688 0 1 45472
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  input64
timestamp 1698431365
transform 1 0 216720 0 1 45472
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_3  input65
timestamp 1698431365
transform 1 0 11088 0 1 45472
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input66
timestamp 1698431365
transform 1 0 15120 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input67
timestamp 1698431365
transform 1 0 19152 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input68
timestamp 1698431365
transform 1 0 23184 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input69
timestamp 1698431365
transform 1 0 28224 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input70
timestamp 1698431365
transform 1 0 32032 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input71
timestamp 1698431365
transform 1 0 35840 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input72
timestamp 1698431365
transform 1 0 39648 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input73
timestamp 1698431365
transform 1 0 43456 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input74
timestamp 1698431365
transform 1 0 79632 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input75
timestamp 1698431365
transform 1 0 83664 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input76
timestamp 1698431365
transform 1 0 123984 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input77
timestamp 1698431365
transform 1 0 128016 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input78
timestamp 1698431365
transform 1 0 132048 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input79
timestamp 1698431365
transform -1 0 136752 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input80
timestamp 1698431365
transform -1 0 140784 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input81
timestamp 1698431365
transform -1 0 144816 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input82
timestamp 1698431365
transform 1 0 87696 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input83
timestamp 1698431365
transform 1 0 91728 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input84
timestamp 1698431365
transform 1 0 95760 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input85
timestamp 1698431365
transform 1 0 100576 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input86
timestamp 1698431365
transform 1 0 104384 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input87
timestamp 1698431365
transform 1 0 108192 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input88
timestamp 1698431365
transform 1 0 112000 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input89
timestamp 1698431365
transform 1 0 115920 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input90
timestamp 1698431365
transform 1 0 119952 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input91
timestamp 1698431365
transform -1 0 7728 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output92 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 31136 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output93
timestamp 1698431365
transform -1 0 32704 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output94
timestamp 1698431365
transform -1 0 35616 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output95
timestamp 1698431365
transform -1 0 38864 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output96
timestamp 1698431365
transform -1 0 42560 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output97
timestamp 1698431365
transform -1 0 44240 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output98
timestamp 1698431365
transform -1 0 46928 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output99
timestamp 1698431365
transform -1 0 50176 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output100
timestamp 1698431365
transform -1 0 52304 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output101
timestamp 1698431365
transform -1 0 6608 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output102
timestamp 1698431365
transform 1 0 51744 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output103
timestamp 1698431365
transform 1 0 54880 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output104
timestamp 1698431365
transform 1 0 57456 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output105
timestamp 1698431365
transform 1 0 59360 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output106
timestamp 1698431365
transform 1 0 62832 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output107
timestamp 1698431365
transform 1 0 66304 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output108
timestamp 1698431365
transform 1 0 68208 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output109
timestamp 1698431365
transform 1 0 70784 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output110
timestamp 1698431365
transform -1 0 76832 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output111
timestamp 1698431365
transform -1 0 79184 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output112
timestamp 1698431365
transform -1 0 81312 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output113
timestamp 1698431365
transform -1 0 84560 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output114
timestamp 1698431365
transform -1 0 87248 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output115
timestamp 1698431365
transform -1 0 88928 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output116
timestamp 1698431365
transform -1 0 152992 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output117
timestamp 1698431365
transform 1 0 152208 0 -1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output118
timestamp 1698431365
transform -1 0 50288 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output119
timestamp 1698431365
transform -1 0 54320 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output120
timestamp 1698431365
transform -1 0 58352 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output121
timestamp 1698431365
transform -1 0 62272 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output122
timestamp 1698431365
transform -1 0 66080 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output123
timestamp 1698431365
transform -1 0 69888 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output124
timestamp 1698431365
transform -1 0 73696 0 1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output125
timestamp 1698431365
transform -1 0 78512 0 -1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_55 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 218624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_56
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 218624 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_57
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 218624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_58
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 218624 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_59
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 218624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_60
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 218624 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_61
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 218624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_62
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 218624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_63
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 218624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_64
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 218624 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_65
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 218624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_66
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 218624 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_67
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 218624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_68
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 218624 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_69
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 218624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_70
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 218624 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_71
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 218624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_72
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 218624 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_73
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 218624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_74
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 218624 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_75
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 218624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_76
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 218624 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_77
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 218624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_78
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 218624 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_79
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 218624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_80
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 218624 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_81
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 218624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_82
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 218624 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_83
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 218624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_84
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 218624 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_85
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 218624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_86
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 218624 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_87
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 218624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_88
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 218624 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_89
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 218624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_90
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 218624 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_91
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 218624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_92
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 218624 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_93
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 218624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_94
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 218624 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_95
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 218624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_96
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 218624 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_97
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 218624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_98
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 218624 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_99
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 218624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_100
timestamp 1698431365
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 218624 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_101
timestamp 1698431365
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 218624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_102
timestamp 1698431365
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 218624 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_103
timestamp 1698431365
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 218624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_104
timestamp 1698431365
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 218624 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_105
timestamp 1698431365
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698431365
transform -1 0 218624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_106
timestamp 1698431365
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698431365
transform -1 0 218624 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_107
timestamp 1698431365
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1698431365
transform -1 0 218624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_108
timestamp 1698431365
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1698431365
transform -1 0 218624 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_109
timestamp 1698431365
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1698431365
transform -1 0 218624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ram_controller_126 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 6832 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ram_controller_127
timestamp 1698431365
transform -1 0 9632 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ram_controller_128
timestamp 1698431365
transform -1 0 12208 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ram_controller_129
timestamp 1698431365
transform -1 0 14896 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ram_controller_130
timestamp 1698431365
transform -1 0 17584 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ram_controller_131
timestamp 1698431365
transform -1 0 20272 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ram_controller_132
timestamp 1698431365
transform -1 0 22960 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ram_controller_133
timestamp 1698431365
transform -1 0 25648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_110 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_111
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_112
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_113
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_114
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_115
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_116
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_117
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_118
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_119
timestamp 1698431365
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_120
timestamp 1698431365
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_121
timestamp 1698431365
transform 1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_122
timestamp 1698431365
transform 1 0 50848 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_123
timestamp 1698431365
transform 1 0 54656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_124
timestamp 1698431365
transform 1 0 58464 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_125
timestamp 1698431365
transform 1 0 62272 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_126
timestamp 1698431365
transform 1 0 66080 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_127
timestamp 1698431365
transform 1 0 69888 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_128
timestamp 1698431365
transform 1 0 73696 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_129
timestamp 1698431365
transform 1 0 77504 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_130
timestamp 1698431365
transform 1 0 81312 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_131
timestamp 1698431365
transform 1 0 85120 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_132
timestamp 1698431365
transform 1 0 88928 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_133
timestamp 1698431365
transform 1 0 92736 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_134
timestamp 1698431365
transform 1 0 96544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_135
timestamp 1698431365
transform 1 0 100352 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_136
timestamp 1698431365
transform 1 0 104160 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_137
timestamp 1698431365
transform 1 0 107968 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_138
timestamp 1698431365
transform 1 0 111776 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_139
timestamp 1698431365
transform 1 0 115584 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_140
timestamp 1698431365
transform 1 0 119392 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_141
timestamp 1698431365
transform 1 0 123200 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_142
timestamp 1698431365
transform 1 0 127008 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_143
timestamp 1698431365
transform 1 0 130816 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_144
timestamp 1698431365
transform 1 0 134624 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_145
timestamp 1698431365
transform 1 0 138432 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_146
timestamp 1698431365
transform 1 0 142240 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_147
timestamp 1698431365
transform 1 0 146048 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_148
timestamp 1698431365
transform 1 0 149856 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_149
timestamp 1698431365
transform 1 0 153664 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_150
timestamp 1698431365
transform 1 0 157472 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_151
timestamp 1698431365
transform 1 0 161280 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_152
timestamp 1698431365
transform 1 0 165088 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_153
timestamp 1698431365
transform 1 0 168896 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_154
timestamp 1698431365
transform 1 0 172704 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_155
timestamp 1698431365
transform 1 0 176512 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_156
timestamp 1698431365
transform 1 0 180320 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_157
timestamp 1698431365
transform 1 0 184128 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_158
timestamp 1698431365
transform 1 0 187936 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_159
timestamp 1698431365
transform 1 0 191744 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_160
timestamp 1698431365
transform 1 0 195552 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_161
timestamp 1698431365
transform 1 0 199360 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_162
timestamp 1698431365
transform 1 0 203168 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_163
timestamp 1698431365
transform 1 0 206976 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_164
timestamp 1698431365
transform 1 0 210784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_165
timestamp 1698431365
transform 1 0 214592 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_166
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_167
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_168
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_169
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_170
timestamp 1698431365
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_171
timestamp 1698431365
transform 1 0 48384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_172
timestamp 1698431365
transform 1 0 56224 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_173
timestamp 1698431365
transform 1 0 64064 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_174
timestamp 1698431365
transform 1 0 71904 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_175
timestamp 1698431365
transform 1 0 79744 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_176
timestamp 1698431365
transform 1 0 87584 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_177
timestamp 1698431365
transform 1 0 95424 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_178
timestamp 1698431365
transform 1 0 103264 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_179
timestamp 1698431365
transform 1 0 111104 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_180
timestamp 1698431365
transform 1 0 118944 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_181
timestamp 1698431365
transform 1 0 126784 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_182
timestamp 1698431365
transform 1 0 134624 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_183
timestamp 1698431365
transform 1 0 142464 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_184
timestamp 1698431365
transform 1 0 150304 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_185
timestamp 1698431365
transform 1 0 158144 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_186
timestamp 1698431365
transform 1 0 165984 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_187
timestamp 1698431365
transform 1 0 173824 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_188
timestamp 1698431365
transform 1 0 181664 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_189
timestamp 1698431365
transform 1 0 189504 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_190
timestamp 1698431365
transform 1 0 197344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_191
timestamp 1698431365
transform 1 0 205184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_192
timestamp 1698431365
transform 1 0 213024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_193
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_194
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_195
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_196
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_197
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_198
timestamp 1698431365
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_199
timestamp 1698431365
transform 1 0 52304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_200
timestamp 1698431365
transform 1 0 60144 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_201
timestamp 1698431365
transform 1 0 67984 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_202
timestamp 1698431365
transform 1 0 75824 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_203
timestamp 1698431365
transform 1 0 83664 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_204
timestamp 1698431365
transform 1 0 91504 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_205
timestamp 1698431365
transform 1 0 99344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_206
timestamp 1698431365
transform 1 0 107184 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_207
timestamp 1698431365
transform 1 0 115024 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_208
timestamp 1698431365
transform 1 0 122864 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_209
timestamp 1698431365
transform 1 0 130704 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_210
timestamp 1698431365
transform 1 0 138544 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_211
timestamp 1698431365
transform 1 0 146384 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_212
timestamp 1698431365
transform 1 0 154224 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_213
timestamp 1698431365
transform 1 0 162064 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_214
timestamp 1698431365
transform 1 0 169904 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_215
timestamp 1698431365
transform 1 0 177744 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_216
timestamp 1698431365
transform 1 0 185584 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_217
timestamp 1698431365
transform 1 0 193424 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_218
timestamp 1698431365
transform 1 0 201264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_219
timestamp 1698431365
transform 1 0 209104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_220
timestamp 1698431365
transform 1 0 216944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_221
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_222
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_223
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_224
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_225
timestamp 1698431365
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_226
timestamp 1698431365
transform 1 0 48384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_227
timestamp 1698431365
transform 1 0 56224 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_228
timestamp 1698431365
transform 1 0 64064 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_229
timestamp 1698431365
transform 1 0 71904 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_230
timestamp 1698431365
transform 1 0 79744 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_231
timestamp 1698431365
transform 1 0 87584 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_232
timestamp 1698431365
transform 1 0 95424 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_233
timestamp 1698431365
transform 1 0 103264 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_234
timestamp 1698431365
transform 1 0 111104 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_235
timestamp 1698431365
transform 1 0 118944 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_236
timestamp 1698431365
transform 1 0 126784 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_237
timestamp 1698431365
transform 1 0 134624 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_238
timestamp 1698431365
transform 1 0 142464 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_239
timestamp 1698431365
transform 1 0 150304 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_240
timestamp 1698431365
transform 1 0 158144 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_241
timestamp 1698431365
transform 1 0 165984 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_242
timestamp 1698431365
transform 1 0 173824 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_243
timestamp 1698431365
transform 1 0 181664 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_244
timestamp 1698431365
transform 1 0 189504 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_245
timestamp 1698431365
transform 1 0 197344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_246
timestamp 1698431365
transform 1 0 205184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_247
timestamp 1698431365
transform 1 0 213024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_248
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_249
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_250
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_251
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_252
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_253
timestamp 1698431365
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_254
timestamp 1698431365
transform 1 0 52304 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_255
timestamp 1698431365
transform 1 0 60144 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_256
timestamp 1698431365
transform 1 0 67984 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_257
timestamp 1698431365
transform 1 0 75824 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_258
timestamp 1698431365
transform 1 0 83664 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_259
timestamp 1698431365
transform 1 0 91504 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_260
timestamp 1698431365
transform 1 0 99344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_261
timestamp 1698431365
transform 1 0 107184 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_262
timestamp 1698431365
transform 1 0 115024 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_263
timestamp 1698431365
transform 1 0 122864 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_264
timestamp 1698431365
transform 1 0 130704 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_265
timestamp 1698431365
transform 1 0 138544 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_266
timestamp 1698431365
transform 1 0 146384 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_267
timestamp 1698431365
transform 1 0 154224 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_268
timestamp 1698431365
transform 1 0 162064 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_269
timestamp 1698431365
transform 1 0 169904 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_270
timestamp 1698431365
transform 1 0 177744 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_271
timestamp 1698431365
transform 1 0 185584 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_272
timestamp 1698431365
transform 1 0 193424 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_273
timestamp 1698431365
transform 1 0 201264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_274
timestamp 1698431365
transform 1 0 209104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_275
timestamp 1698431365
transform 1 0 216944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_276
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_277
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_278
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_279
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_280
timestamp 1698431365
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_281
timestamp 1698431365
transform 1 0 48384 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_282
timestamp 1698431365
transform 1 0 56224 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_283
timestamp 1698431365
transform 1 0 64064 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_284
timestamp 1698431365
transform 1 0 71904 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_285
timestamp 1698431365
transform 1 0 79744 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_286
timestamp 1698431365
transform 1 0 87584 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_287
timestamp 1698431365
transform 1 0 95424 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_288
timestamp 1698431365
transform 1 0 103264 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_289
timestamp 1698431365
transform 1 0 111104 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_290
timestamp 1698431365
transform 1 0 118944 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_291
timestamp 1698431365
transform 1 0 126784 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_292
timestamp 1698431365
transform 1 0 134624 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_293
timestamp 1698431365
transform 1 0 142464 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_294
timestamp 1698431365
transform 1 0 150304 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_295
timestamp 1698431365
transform 1 0 158144 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_296
timestamp 1698431365
transform 1 0 165984 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_297
timestamp 1698431365
transform 1 0 173824 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_298
timestamp 1698431365
transform 1 0 181664 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_299
timestamp 1698431365
transform 1 0 189504 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_300
timestamp 1698431365
transform 1 0 197344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_301
timestamp 1698431365
transform 1 0 205184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_302
timestamp 1698431365
transform 1 0 213024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_303
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_304
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_305
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_306
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_307
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_308
timestamp 1698431365
transform 1 0 44464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_309
timestamp 1698431365
transform 1 0 52304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_310
timestamp 1698431365
transform 1 0 60144 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_311
timestamp 1698431365
transform 1 0 67984 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_312
timestamp 1698431365
transform 1 0 75824 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_313
timestamp 1698431365
transform 1 0 83664 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_314
timestamp 1698431365
transform 1 0 91504 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_315
timestamp 1698431365
transform 1 0 99344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_316
timestamp 1698431365
transform 1 0 107184 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_317
timestamp 1698431365
transform 1 0 115024 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_318
timestamp 1698431365
transform 1 0 122864 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_319
timestamp 1698431365
transform 1 0 130704 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_320
timestamp 1698431365
transform 1 0 138544 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_321
timestamp 1698431365
transform 1 0 146384 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_322
timestamp 1698431365
transform 1 0 154224 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_323
timestamp 1698431365
transform 1 0 162064 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_324
timestamp 1698431365
transform 1 0 169904 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_325
timestamp 1698431365
transform 1 0 177744 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_326
timestamp 1698431365
transform 1 0 185584 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_327
timestamp 1698431365
transform 1 0 193424 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_328
timestamp 1698431365
transform 1 0 201264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_329
timestamp 1698431365
transform 1 0 209104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_330
timestamp 1698431365
transform 1 0 216944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_331
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_332
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_333
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_334
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_335
timestamp 1698431365
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_336
timestamp 1698431365
transform 1 0 48384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_337
timestamp 1698431365
transform 1 0 56224 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_338
timestamp 1698431365
transform 1 0 64064 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_339
timestamp 1698431365
transform 1 0 71904 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_340
timestamp 1698431365
transform 1 0 79744 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_341
timestamp 1698431365
transform 1 0 87584 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_342
timestamp 1698431365
transform 1 0 95424 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_343
timestamp 1698431365
transform 1 0 103264 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_344
timestamp 1698431365
transform 1 0 111104 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_345
timestamp 1698431365
transform 1 0 118944 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_346
timestamp 1698431365
transform 1 0 126784 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_347
timestamp 1698431365
transform 1 0 134624 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_348
timestamp 1698431365
transform 1 0 142464 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_349
timestamp 1698431365
transform 1 0 150304 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_350
timestamp 1698431365
transform 1 0 158144 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_351
timestamp 1698431365
transform 1 0 165984 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_352
timestamp 1698431365
transform 1 0 173824 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_353
timestamp 1698431365
transform 1 0 181664 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_354
timestamp 1698431365
transform 1 0 189504 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_355
timestamp 1698431365
transform 1 0 197344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_356
timestamp 1698431365
transform 1 0 205184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_357
timestamp 1698431365
transform 1 0 213024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_358
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_359
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_360
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_361
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_362
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_363
timestamp 1698431365
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_364
timestamp 1698431365
transform 1 0 52304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_365
timestamp 1698431365
transform 1 0 60144 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_366
timestamp 1698431365
transform 1 0 67984 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_367
timestamp 1698431365
transform 1 0 75824 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_368
timestamp 1698431365
transform 1 0 83664 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_369
timestamp 1698431365
transform 1 0 91504 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_370
timestamp 1698431365
transform 1 0 99344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_371
timestamp 1698431365
transform 1 0 107184 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_372
timestamp 1698431365
transform 1 0 115024 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_373
timestamp 1698431365
transform 1 0 122864 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_374
timestamp 1698431365
transform 1 0 130704 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_375
timestamp 1698431365
transform 1 0 138544 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_376
timestamp 1698431365
transform 1 0 146384 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_377
timestamp 1698431365
transform 1 0 154224 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_378
timestamp 1698431365
transform 1 0 162064 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_379
timestamp 1698431365
transform 1 0 169904 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_380
timestamp 1698431365
transform 1 0 177744 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_381
timestamp 1698431365
transform 1 0 185584 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_382
timestamp 1698431365
transform 1 0 193424 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_383
timestamp 1698431365
transform 1 0 201264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_384
timestamp 1698431365
transform 1 0 209104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_385
timestamp 1698431365
transform 1 0 216944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_386
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_387
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_388
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_389
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_390
timestamp 1698431365
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_391
timestamp 1698431365
transform 1 0 48384 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_392
timestamp 1698431365
transform 1 0 56224 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_393
timestamp 1698431365
transform 1 0 64064 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_394
timestamp 1698431365
transform 1 0 71904 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_395
timestamp 1698431365
transform 1 0 79744 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_396
timestamp 1698431365
transform 1 0 87584 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_397
timestamp 1698431365
transform 1 0 95424 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_398
timestamp 1698431365
transform 1 0 103264 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_399
timestamp 1698431365
transform 1 0 111104 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_400
timestamp 1698431365
transform 1 0 118944 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_401
timestamp 1698431365
transform 1 0 126784 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_402
timestamp 1698431365
transform 1 0 134624 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_403
timestamp 1698431365
transform 1 0 142464 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_404
timestamp 1698431365
transform 1 0 150304 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_405
timestamp 1698431365
transform 1 0 158144 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_406
timestamp 1698431365
transform 1 0 165984 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_407
timestamp 1698431365
transform 1 0 173824 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_408
timestamp 1698431365
transform 1 0 181664 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_409
timestamp 1698431365
transform 1 0 189504 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_410
timestamp 1698431365
transform 1 0 197344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_411
timestamp 1698431365
transform 1 0 205184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_412
timestamp 1698431365
transform 1 0 213024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_413
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_414
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_415
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_416
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_417
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_418
timestamp 1698431365
transform 1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_419
timestamp 1698431365
transform 1 0 52304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_420
timestamp 1698431365
transform 1 0 60144 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_421
timestamp 1698431365
transform 1 0 67984 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_422
timestamp 1698431365
transform 1 0 75824 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_423
timestamp 1698431365
transform 1 0 83664 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_424
timestamp 1698431365
transform 1 0 91504 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_425
timestamp 1698431365
transform 1 0 99344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_426
timestamp 1698431365
transform 1 0 107184 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_427
timestamp 1698431365
transform 1 0 115024 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_428
timestamp 1698431365
transform 1 0 122864 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_429
timestamp 1698431365
transform 1 0 130704 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_430
timestamp 1698431365
transform 1 0 138544 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_431
timestamp 1698431365
transform 1 0 146384 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_432
timestamp 1698431365
transform 1 0 154224 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_433
timestamp 1698431365
transform 1 0 162064 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_434
timestamp 1698431365
transform 1 0 169904 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_435
timestamp 1698431365
transform 1 0 177744 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_436
timestamp 1698431365
transform 1 0 185584 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_437
timestamp 1698431365
transform 1 0 193424 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_438
timestamp 1698431365
transform 1 0 201264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_439
timestamp 1698431365
transform 1 0 209104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_440
timestamp 1698431365
transform 1 0 216944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_441
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_442
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_443
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_444
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_445
timestamp 1698431365
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_446
timestamp 1698431365
transform 1 0 48384 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_447
timestamp 1698431365
transform 1 0 56224 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_448
timestamp 1698431365
transform 1 0 64064 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_449
timestamp 1698431365
transform 1 0 71904 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_450
timestamp 1698431365
transform 1 0 79744 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_451
timestamp 1698431365
transform 1 0 87584 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_452
timestamp 1698431365
transform 1 0 95424 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_453
timestamp 1698431365
transform 1 0 103264 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_454
timestamp 1698431365
transform 1 0 111104 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_455
timestamp 1698431365
transform 1 0 118944 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_456
timestamp 1698431365
transform 1 0 126784 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_457
timestamp 1698431365
transform 1 0 134624 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_458
timestamp 1698431365
transform 1 0 142464 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_459
timestamp 1698431365
transform 1 0 150304 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_460
timestamp 1698431365
transform 1 0 158144 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_461
timestamp 1698431365
transform 1 0 165984 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_462
timestamp 1698431365
transform 1 0 173824 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_463
timestamp 1698431365
transform 1 0 181664 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_464
timestamp 1698431365
transform 1 0 189504 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_465
timestamp 1698431365
transform 1 0 197344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_466
timestamp 1698431365
transform 1 0 205184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_467
timestamp 1698431365
transform 1 0 213024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_468
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_469
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_470
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_471
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_472
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_473
timestamp 1698431365
transform 1 0 44464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_474
timestamp 1698431365
transform 1 0 52304 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_475
timestamp 1698431365
transform 1 0 60144 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_476
timestamp 1698431365
transform 1 0 67984 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_477
timestamp 1698431365
transform 1 0 75824 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_478
timestamp 1698431365
transform 1 0 83664 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_479
timestamp 1698431365
transform 1 0 91504 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_480
timestamp 1698431365
transform 1 0 99344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_481
timestamp 1698431365
transform 1 0 107184 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_482
timestamp 1698431365
transform 1 0 115024 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_483
timestamp 1698431365
transform 1 0 122864 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_484
timestamp 1698431365
transform 1 0 130704 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_485
timestamp 1698431365
transform 1 0 138544 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_486
timestamp 1698431365
transform 1 0 146384 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_487
timestamp 1698431365
transform 1 0 154224 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_488
timestamp 1698431365
transform 1 0 162064 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_489
timestamp 1698431365
transform 1 0 169904 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_490
timestamp 1698431365
transform 1 0 177744 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_491
timestamp 1698431365
transform 1 0 185584 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_492
timestamp 1698431365
transform 1 0 193424 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_493
timestamp 1698431365
transform 1 0 201264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_494
timestamp 1698431365
transform 1 0 209104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_495
timestamp 1698431365
transform 1 0 216944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_496
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_497
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_498
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_499
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_500
timestamp 1698431365
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_501
timestamp 1698431365
transform 1 0 48384 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_502
timestamp 1698431365
transform 1 0 56224 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_503
timestamp 1698431365
transform 1 0 64064 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_504
timestamp 1698431365
transform 1 0 71904 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_505
timestamp 1698431365
transform 1 0 79744 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_506
timestamp 1698431365
transform 1 0 87584 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_507
timestamp 1698431365
transform 1 0 95424 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_508
timestamp 1698431365
transform 1 0 103264 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_509
timestamp 1698431365
transform 1 0 111104 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_510
timestamp 1698431365
transform 1 0 118944 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_511
timestamp 1698431365
transform 1 0 126784 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_512
timestamp 1698431365
transform 1 0 134624 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_513
timestamp 1698431365
transform 1 0 142464 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_514
timestamp 1698431365
transform 1 0 150304 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_515
timestamp 1698431365
transform 1 0 158144 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_516
timestamp 1698431365
transform 1 0 165984 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_517
timestamp 1698431365
transform 1 0 173824 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_518
timestamp 1698431365
transform 1 0 181664 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_519
timestamp 1698431365
transform 1 0 189504 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_520
timestamp 1698431365
transform 1 0 197344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_521
timestamp 1698431365
transform 1 0 205184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_522
timestamp 1698431365
transform 1 0 213024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_523
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_524
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_525
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_526
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_527
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_528
timestamp 1698431365
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_529
timestamp 1698431365
transform 1 0 52304 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_530
timestamp 1698431365
transform 1 0 60144 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_531
timestamp 1698431365
transform 1 0 67984 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_532
timestamp 1698431365
transform 1 0 75824 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_533
timestamp 1698431365
transform 1 0 83664 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_534
timestamp 1698431365
transform 1 0 91504 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_535
timestamp 1698431365
transform 1 0 99344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_536
timestamp 1698431365
transform 1 0 107184 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_537
timestamp 1698431365
transform 1 0 115024 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_538
timestamp 1698431365
transform 1 0 122864 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_539
timestamp 1698431365
transform 1 0 130704 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_540
timestamp 1698431365
transform 1 0 138544 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_541
timestamp 1698431365
transform 1 0 146384 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_542
timestamp 1698431365
transform 1 0 154224 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_543
timestamp 1698431365
transform 1 0 162064 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_544
timestamp 1698431365
transform 1 0 169904 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_545
timestamp 1698431365
transform 1 0 177744 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_546
timestamp 1698431365
transform 1 0 185584 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_547
timestamp 1698431365
transform 1 0 193424 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_548
timestamp 1698431365
transform 1 0 201264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_549
timestamp 1698431365
transform 1 0 209104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_550
timestamp 1698431365
transform 1 0 216944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_551
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_552
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_553
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_554
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_555
timestamp 1698431365
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_556
timestamp 1698431365
transform 1 0 48384 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_557
timestamp 1698431365
transform 1 0 56224 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_558
timestamp 1698431365
transform 1 0 64064 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_559
timestamp 1698431365
transform 1 0 71904 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_560
timestamp 1698431365
transform 1 0 79744 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_561
timestamp 1698431365
transform 1 0 87584 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_562
timestamp 1698431365
transform 1 0 95424 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_563
timestamp 1698431365
transform 1 0 103264 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_564
timestamp 1698431365
transform 1 0 111104 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_565
timestamp 1698431365
transform 1 0 118944 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_566
timestamp 1698431365
transform 1 0 126784 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_567
timestamp 1698431365
transform 1 0 134624 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_568
timestamp 1698431365
transform 1 0 142464 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_569
timestamp 1698431365
transform 1 0 150304 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_570
timestamp 1698431365
transform 1 0 158144 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_571
timestamp 1698431365
transform 1 0 165984 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_572
timestamp 1698431365
transform 1 0 173824 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_573
timestamp 1698431365
transform 1 0 181664 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_574
timestamp 1698431365
transform 1 0 189504 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_575
timestamp 1698431365
transform 1 0 197344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_576
timestamp 1698431365
transform 1 0 205184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_577
timestamp 1698431365
transform 1 0 213024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_578
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_579
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_580
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_581
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_582
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_583
timestamp 1698431365
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_584
timestamp 1698431365
transform 1 0 52304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_585
timestamp 1698431365
transform 1 0 60144 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_586
timestamp 1698431365
transform 1 0 67984 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_587
timestamp 1698431365
transform 1 0 75824 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_588
timestamp 1698431365
transform 1 0 83664 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_589
timestamp 1698431365
transform 1 0 91504 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_590
timestamp 1698431365
transform 1 0 99344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_591
timestamp 1698431365
transform 1 0 107184 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_592
timestamp 1698431365
transform 1 0 115024 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_593
timestamp 1698431365
transform 1 0 122864 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_594
timestamp 1698431365
transform 1 0 130704 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_595
timestamp 1698431365
transform 1 0 138544 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_596
timestamp 1698431365
transform 1 0 146384 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_597
timestamp 1698431365
transform 1 0 154224 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_598
timestamp 1698431365
transform 1 0 162064 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_599
timestamp 1698431365
transform 1 0 169904 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_600
timestamp 1698431365
transform 1 0 177744 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_601
timestamp 1698431365
transform 1 0 185584 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_602
timestamp 1698431365
transform 1 0 193424 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_603
timestamp 1698431365
transform 1 0 201264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_604
timestamp 1698431365
transform 1 0 209104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_605
timestamp 1698431365
transform 1 0 216944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_606
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_607
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_608
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_609
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_610
timestamp 1698431365
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_611
timestamp 1698431365
transform 1 0 48384 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_612
timestamp 1698431365
transform 1 0 56224 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_613
timestamp 1698431365
transform 1 0 64064 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_614
timestamp 1698431365
transform 1 0 71904 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_615
timestamp 1698431365
transform 1 0 79744 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_616
timestamp 1698431365
transform 1 0 87584 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_617
timestamp 1698431365
transform 1 0 95424 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_618
timestamp 1698431365
transform 1 0 103264 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_619
timestamp 1698431365
transform 1 0 111104 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_620
timestamp 1698431365
transform 1 0 118944 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_621
timestamp 1698431365
transform 1 0 126784 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_622
timestamp 1698431365
transform 1 0 134624 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_623
timestamp 1698431365
transform 1 0 142464 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_624
timestamp 1698431365
transform 1 0 150304 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_625
timestamp 1698431365
transform 1 0 158144 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_626
timestamp 1698431365
transform 1 0 165984 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_627
timestamp 1698431365
transform 1 0 173824 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_628
timestamp 1698431365
transform 1 0 181664 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_629
timestamp 1698431365
transform 1 0 189504 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_630
timestamp 1698431365
transform 1 0 197344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_631
timestamp 1698431365
transform 1 0 205184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_632
timestamp 1698431365
transform 1 0 213024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_633
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_634
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_635
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_636
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_637
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_638
timestamp 1698431365
transform 1 0 44464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_639
timestamp 1698431365
transform 1 0 52304 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_640
timestamp 1698431365
transform 1 0 60144 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_641
timestamp 1698431365
transform 1 0 67984 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_642
timestamp 1698431365
transform 1 0 75824 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_643
timestamp 1698431365
transform 1 0 83664 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_644
timestamp 1698431365
transform 1 0 91504 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_645
timestamp 1698431365
transform 1 0 99344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_646
timestamp 1698431365
transform 1 0 107184 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_647
timestamp 1698431365
transform 1 0 115024 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_648
timestamp 1698431365
transform 1 0 122864 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_649
timestamp 1698431365
transform 1 0 130704 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_650
timestamp 1698431365
transform 1 0 138544 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_651
timestamp 1698431365
transform 1 0 146384 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_652
timestamp 1698431365
transform 1 0 154224 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_653
timestamp 1698431365
transform 1 0 162064 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_654
timestamp 1698431365
transform 1 0 169904 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_655
timestamp 1698431365
transform 1 0 177744 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_656
timestamp 1698431365
transform 1 0 185584 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_657
timestamp 1698431365
transform 1 0 193424 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_658
timestamp 1698431365
transform 1 0 201264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_659
timestamp 1698431365
transform 1 0 209104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_660
timestamp 1698431365
transform 1 0 216944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_661
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_662
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_663
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_664
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_665
timestamp 1698431365
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_666
timestamp 1698431365
transform 1 0 48384 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_667
timestamp 1698431365
transform 1 0 56224 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_668
timestamp 1698431365
transform 1 0 64064 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_669
timestamp 1698431365
transform 1 0 71904 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_670
timestamp 1698431365
transform 1 0 79744 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_671
timestamp 1698431365
transform 1 0 87584 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_672
timestamp 1698431365
transform 1 0 95424 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_673
timestamp 1698431365
transform 1 0 103264 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_674
timestamp 1698431365
transform 1 0 111104 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_675
timestamp 1698431365
transform 1 0 118944 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_676
timestamp 1698431365
transform 1 0 126784 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_677
timestamp 1698431365
transform 1 0 134624 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_678
timestamp 1698431365
transform 1 0 142464 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_679
timestamp 1698431365
transform 1 0 150304 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_680
timestamp 1698431365
transform 1 0 158144 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_681
timestamp 1698431365
transform 1 0 165984 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_682
timestamp 1698431365
transform 1 0 173824 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_683
timestamp 1698431365
transform 1 0 181664 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_684
timestamp 1698431365
transform 1 0 189504 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_685
timestamp 1698431365
transform 1 0 197344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_686
timestamp 1698431365
transform 1 0 205184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_687
timestamp 1698431365
transform 1 0 213024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_688
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_689
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_690
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_691
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_692
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_693
timestamp 1698431365
transform 1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_694
timestamp 1698431365
transform 1 0 52304 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_695
timestamp 1698431365
transform 1 0 60144 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_696
timestamp 1698431365
transform 1 0 67984 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_697
timestamp 1698431365
transform 1 0 75824 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_698
timestamp 1698431365
transform 1 0 83664 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_699
timestamp 1698431365
transform 1 0 91504 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_700
timestamp 1698431365
transform 1 0 99344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_701
timestamp 1698431365
transform 1 0 107184 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_702
timestamp 1698431365
transform 1 0 115024 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_703
timestamp 1698431365
transform 1 0 122864 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_704
timestamp 1698431365
transform 1 0 130704 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_705
timestamp 1698431365
transform 1 0 138544 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_706
timestamp 1698431365
transform 1 0 146384 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_707
timestamp 1698431365
transform 1 0 154224 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_708
timestamp 1698431365
transform 1 0 162064 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_709
timestamp 1698431365
transform 1 0 169904 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_710
timestamp 1698431365
transform 1 0 177744 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_711
timestamp 1698431365
transform 1 0 185584 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_712
timestamp 1698431365
transform 1 0 193424 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_713
timestamp 1698431365
transform 1 0 201264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_714
timestamp 1698431365
transform 1 0 209104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_715
timestamp 1698431365
transform 1 0 216944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_716
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_717
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_718
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_719
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_720
timestamp 1698431365
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_721
timestamp 1698431365
transform 1 0 48384 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_722
timestamp 1698431365
transform 1 0 56224 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_723
timestamp 1698431365
transform 1 0 64064 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_724
timestamp 1698431365
transform 1 0 71904 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_725
timestamp 1698431365
transform 1 0 79744 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_726
timestamp 1698431365
transform 1 0 87584 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_727
timestamp 1698431365
transform 1 0 95424 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_728
timestamp 1698431365
transform 1 0 103264 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_729
timestamp 1698431365
transform 1 0 111104 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_730
timestamp 1698431365
transform 1 0 118944 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_731
timestamp 1698431365
transform 1 0 126784 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_732
timestamp 1698431365
transform 1 0 134624 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_733
timestamp 1698431365
transform 1 0 142464 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_734
timestamp 1698431365
transform 1 0 150304 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_735
timestamp 1698431365
transform 1 0 158144 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_736
timestamp 1698431365
transform 1 0 165984 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_737
timestamp 1698431365
transform 1 0 173824 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_738
timestamp 1698431365
transform 1 0 181664 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_739
timestamp 1698431365
transform 1 0 189504 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_740
timestamp 1698431365
transform 1 0 197344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_741
timestamp 1698431365
transform 1 0 205184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_742
timestamp 1698431365
transform 1 0 213024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_743
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_744
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_745
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_746
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_747
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_748
timestamp 1698431365
transform 1 0 44464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_749
timestamp 1698431365
transform 1 0 52304 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_750
timestamp 1698431365
transform 1 0 60144 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_751
timestamp 1698431365
transform 1 0 67984 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_752
timestamp 1698431365
transform 1 0 75824 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_753
timestamp 1698431365
transform 1 0 83664 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_754
timestamp 1698431365
transform 1 0 91504 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_755
timestamp 1698431365
transform 1 0 99344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_756
timestamp 1698431365
transform 1 0 107184 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_757
timestamp 1698431365
transform 1 0 115024 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_758
timestamp 1698431365
transform 1 0 122864 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_759
timestamp 1698431365
transform 1 0 130704 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_760
timestamp 1698431365
transform 1 0 138544 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_761
timestamp 1698431365
transform 1 0 146384 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_762
timestamp 1698431365
transform 1 0 154224 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_763
timestamp 1698431365
transform 1 0 162064 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_764
timestamp 1698431365
transform 1 0 169904 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_765
timestamp 1698431365
transform 1 0 177744 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_766
timestamp 1698431365
transform 1 0 185584 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_767
timestamp 1698431365
transform 1 0 193424 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_768
timestamp 1698431365
transform 1 0 201264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_769
timestamp 1698431365
transform 1 0 209104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_770
timestamp 1698431365
transform 1 0 216944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_771
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_772
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_773
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_774
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_775
timestamp 1698431365
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_776
timestamp 1698431365
transform 1 0 48384 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_777
timestamp 1698431365
transform 1 0 56224 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_778
timestamp 1698431365
transform 1 0 64064 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_779
timestamp 1698431365
transform 1 0 71904 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_780
timestamp 1698431365
transform 1 0 79744 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_781
timestamp 1698431365
transform 1 0 87584 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_782
timestamp 1698431365
transform 1 0 95424 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_783
timestamp 1698431365
transform 1 0 103264 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_784
timestamp 1698431365
transform 1 0 111104 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_785
timestamp 1698431365
transform 1 0 118944 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_786
timestamp 1698431365
transform 1 0 126784 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_787
timestamp 1698431365
transform 1 0 134624 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_788
timestamp 1698431365
transform 1 0 142464 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_789
timestamp 1698431365
transform 1 0 150304 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_790
timestamp 1698431365
transform 1 0 158144 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_791
timestamp 1698431365
transform 1 0 165984 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_792
timestamp 1698431365
transform 1 0 173824 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_793
timestamp 1698431365
transform 1 0 181664 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_794
timestamp 1698431365
transform 1 0 189504 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_795
timestamp 1698431365
transform 1 0 197344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_796
timestamp 1698431365
transform 1 0 205184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_797
timestamp 1698431365
transform 1 0 213024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_798
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_799
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_800
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_801
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_802
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_803
timestamp 1698431365
transform 1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_804
timestamp 1698431365
transform 1 0 52304 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_805
timestamp 1698431365
transform 1 0 60144 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_806
timestamp 1698431365
transform 1 0 67984 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_807
timestamp 1698431365
transform 1 0 75824 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_808
timestamp 1698431365
transform 1 0 83664 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_809
timestamp 1698431365
transform 1 0 91504 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_810
timestamp 1698431365
transform 1 0 99344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_811
timestamp 1698431365
transform 1 0 107184 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_812
timestamp 1698431365
transform 1 0 115024 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_813
timestamp 1698431365
transform 1 0 122864 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_814
timestamp 1698431365
transform 1 0 130704 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_815
timestamp 1698431365
transform 1 0 138544 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_816
timestamp 1698431365
transform 1 0 146384 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_817
timestamp 1698431365
transform 1 0 154224 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_818
timestamp 1698431365
transform 1 0 162064 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_819
timestamp 1698431365
transform 1 0 169904 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_820
timestamp 1698431365
transform 1 0 177744 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_821
timestamp 1698431365
transform 1 0 185584 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_822
timestamp 1698431365
transform 1 0 193424 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_823
timestamp 1698431365
transform 1 0 201264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_824
timestamp 1698431365
transform 1 0 209104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_825
timestamp 1698431365
transform 1 0 216944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_826
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_827
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_828
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_829
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_830
timestamp 1698431365
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_831
timestamp 1698431365
transform 1 0 48384 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_832
timestamp 1698431365
transform 1 0 56224 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_833
timestamp 1698431365
transform 1 0 64064 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_834
timestamp 1698431365
transform 1 0 71904 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_835
timestamp 1698431365
transform 1 0 79744 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_836
timestamp 1698431365
transform 1 0 87584 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_837
timestamp 1698431365
transform 1 0 95424 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_838
timestamp 1698431365
transform 1 0 103264 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_839
timestamp 1698431365
transform 1 0 111104 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_840
timestamp 1698431365
transform 1 0 118944 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_841
timestamp 1698431365
transform 1 0 126784 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_842
timestamp 1698431365
transform 1 0 134624 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_843
timestamp 1698431365
transform 1 0 142464 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_844
timestamp 1698431365
transform 1 0 150304 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_845
timestamp 1698431365
transform 1 0 158144 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_846
timestamp 1698431365
transform 1 0 165984 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_847
timestamp 1698431365
transform 1 0 173824 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_848
timestamp 1698431365
transform 1 0 181664 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_849
timestamp 1698431365
transform 1 0 189504 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_850
timestamp 1698431365
transform 1 0 197344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_851
timestamp 1698431365
transform 1 0 205184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_852
timestamp 1698431365
transform 1 0 213024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_853
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_854
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_855
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_856
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_857
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_858
timestamp 1698431365
transform 1 0 44464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_859
timestamp 1698431365
transform 1 0 52304 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_860
timestamp 1698431365
transform 1 0 60144 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_861
timestamp 1698431365
transform 1 0 67984 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_862
timestamp 1698431365
transform 1 0 75824 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_863
timestamp 1698431365
transform 1 0 83664 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_864
timestamp 1698431365
transform 1 0 91504 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_865
timestamp 1698431365
transform 1 0 99344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_866
timestamp 1698431365
transform 1 0 107184 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_867
timestamp 1698431365
transform 1 0 115024 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_868
timestamp 1698431365
transform 1 0 122864 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_869
timestamp 1698431365
transform 1 0 130704 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_870
timestamp 1698431365
transform 1 0 138544 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_871
timestamp 1698431365
transform 1 0 146384 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_872
timestamp 1698431365
transform 1 0 154224 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_873
timestamp 1698431365
transform 1 0 162064 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_874
timestamp 1698431365
transform 1 0 169904 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_875
timestamp 1698431365
transform 1 0 177744 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_876
timestamp 1698431365
transform 1 0 185584 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_877
timestamp 1698431365
transform 1 0 193424 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_878
timestamp 1698431365
transform 1 0 201264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_879
timestamp 1698431365
transform 1 0 209104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_880
timestamp 1698431365
transform 1 0 216944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_881
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_882
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_883
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_884
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_885
timestamp 1698431365
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_886
timestamp 1698431365
transform 1 0 48384 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_887
timestamp 1698431365
transform 1 0 56224 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_888
timestamp 1698431365
transform 1 0 64064 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_889
timestamp 1698431365
transform 1 0 71904 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_890
timestamp 1698431365
transform 1 0 79744 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_891
timestamp 1698431365
transform 1 0 87584 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_892
timestamp 1698431365
transform 1 0 95424 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_893
timestamp 1698431365
transform 1 0 103264 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_894
timestamp 1698431365
transform 1 0 111104 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_895
timestamp 1698431365
transform 1 0 118944 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_896
timestamp 1698431365
transform 1 0 126784 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_897
timestamp 1698431365
transform 1 0 134624 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_898
timestamp 1698431365
transform 1 0 142464 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_899
timestamp 1698431365
transform 1 0 150304 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_900
timestamp 1698431365
transform 1 0 158144 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_901
timestamp 1698431365
transform 1 0 165984 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_902
timestamp 1698431365
transform 1 0 173824 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_903
timestamp 1698431365
transform 1 0 181664 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_904
timestamp 1698431365
transform 1 0 189504 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_905
timestamp 1698431365
transform 1 0 197344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_906
timestamp 1698431365
transform 1 0 205184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_907
timestamp 1698431365
transform 1 0 213024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_908
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_909
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_910
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_911
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_912
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_913
timestamp 1698431365
transform 1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_914
timestamp 1698431365
transform 1 0 52304 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_915
timestamp 1698431365
transform 1 0 60144 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_916
timestamp 1698431365
transform 1 0 67984 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_917
timestamp 1698431365
transform 1 0 75824 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_918
timestamp 1698431365
transform 1 0 83664 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_919
timestamp 1698431365
transform 1 0 91504 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_920
timestamp 1698431365
transform 1 0 99344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_921
timestamp 1698431365
transform 1 0 107184 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_922
timestamp 1698431365
transform 1 0 115024 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_923
timestamp 1698431365
transform 1 0 122864 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_924
timestamp 1698431365
transform 1 0 130704 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_925
timestamp 1698431365
transform 1 0 138544 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_926
timestamp 1698431365
transform 1 0 146384 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_927
timestamp 1698431365
transform 1 0 154224 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_928
timestamp 1698431365
transform 1 0 162064 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_929
timestamp 1698431365
transform 1 0 169904 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_930
timestamp 1698431365
transform 1 0 177744 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_931
timestamp 1698431365
transform 1 0 185584 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_932
timestamp 1698431365
transform 1 0 193424 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_933
timestamp 1698431365
transform 1 0 201264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_934
timestamp 1698431365
transform 1 0 209104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_935
timestamp 1698431365
transform 1 0 216944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_936
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_937
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_938
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_939
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_940
timestamp 1698431365
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_941
timestamp 1698431365
transform 1 0 48384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_942
timestamp 1698431365
transform 1 0 56224 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_943
timestamp 1698431365
transform 1 0 64064 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_944
timestamp 1698431365
transform 1 0 71904 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_945
timestamp 1698431365
transform 1 0 79744 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_946
timestamp 1698431365
transform 1 0 87584 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_947
timestamp 1698431365
transform 1 0 95424 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_948
timestamp 1698431365
transform 1 0 103264 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_949
timestamp 1698431365
transform 1 0 111104 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_950
timestamp 1698431365
transform 1 0 118944 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_951
timestamp 1698431365
transform 1 0 126784 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_952
timestamp 1698431365
transform 1 0 134624 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_953
timestamp 1698431365
transform 1 0 142464 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_954
timestamp 1698431365
transform 1 0 150304 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_955
timestamp 1698431365
transform 1 0 158144 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_956
timestamp 1698431365
transform 1 0 165984 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_957
timestamp 1698431365
transform 1 0 173824 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_958
timestamp 1698431365
transform 1 0 181664 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_959
timestamp 1698431365
transform 1 0 189504 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_960
timestamp 1698431365
transform 1 0 197344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_961
timestamp 1698431365
transform 1 0 205184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_962
timestamp 1698431365
transform 1 0 213024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_963
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_964
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_965
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_966
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_967
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_968
timestamp 1698431365
transform 1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_969
timestamp 1698431365
transform 1 0 52304 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_970
timestamp 1698431365
transform 1 0 60144 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_971
timestamp 1698431365
transform 1 0 67984 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_972
timestamp 1698431365
transform 1 0 75824 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_973
timestamp 1698431365
transform 1 0 83664 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_974
timestamp 1698431365
transform 1 0 91504 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_975
timestamp 1698431365
transform 1 0 99344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_976
timestamp 1698431365
transform 1 0 107184 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_977
timestamp 1698431365
transform 1 0 115024 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_978
timestamp 1698431365
transform 1 0 122864 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_979
timestamp 1698431365
transform 1 0 130704 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_980
timestamp 1698431365
transform 1 0 138544 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_981
timestamp 1698431365
transform 1 0 146384 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_982
timestamp 1698431365
transform 1 0 154224 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_983
timestamp 1698431365
transform 1 0 162064 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_984
timestamp 1698431365
transform 1 0 169904 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_985
timestamp 1698431365
transform 1 0 177744 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_986
timestamp 1698431365
transform 1 0 185584 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_987
timestamp 1698431365
transform 1 0 193424 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_988
timestamp 1698431365
transform 1 0 201264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_989
timestamp 1698431365
transform 1 0 209104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_990
timestamp 1698431365
transform 1 0 216944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_991
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_992
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_993
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_994
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_995
timestamp 1698431365
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_996
timestamp 1698431365
transform 1 0 48384 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_997
timestamp 1698431365
transform 1 0 56224 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_998
timestamp 1698431365
transform 1 0 64064 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_999
timestamp 1698431365
transform 1 0 71904 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1000
timestamp 1698431365
transform 1 0 79744 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1001
timestamp 1698431365
transform 1 0 87584 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1002
timestamp 1698431365
transform 1 0 95424 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1003
timestamp 1698431365
transform 1 0 103264 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1004
timestamp 1698431365
transform 1 0 111104 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1005
timestamp 1698431365
transform 1 0 118944 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1006
timestamp 1698431365
transform 1 0 126784 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1007
timestamp 1698431365
transform 1 0 134624 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1008
timestamp 1698431365
transform 1 0 142464 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1009
timestamp 1698431365
transform 1 0 150304 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1010
timestamp 1698431365
transform 1 0 158144 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1011
timestamp 1698431365
transform 1 0 165984 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1012
timestamp 1698431365
transform 1 0 173824 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1013
timestamp 1698431365
transform 1 0 181664 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1014
timestamp 1698431365
transform 1 0 189504 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1015
timestamp 1698431365
transform 1 0 197344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1016
timestamp 1698431365
transform 1 0 205184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_1017
timestamp 1698431365
transform 1 0 213024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1018
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1019
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1020
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1021
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1022
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1023
timestamp 1698431365
transform 1 0 44464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1024
timestamp 1698431365
transform 1 0 52304 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1025
timestamp 1698431365
transform 1 0 60144 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1026
timestamp 1698431365
transform 1 0 67984 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1027
timestamp 1698431365
transform 1 0 75824 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1028
timestamp 1698431365
transform 1 0 83664 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1029
timestamp 1698431365
transform 1 0 91504 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1030
timestamp 1698431365
transform 1 0 99344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1031
timestamp 1698431365
transform 1 0 107184 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1032
timestamp 1698431365
transform 1 0 115024 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1033
timestamp 1698431365
transform 1 0 122864 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1034
timestamp 1698431365
transform 1 0 130704 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1035
timestamp 1698431365
transform 1 0 138544 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1036
timestamp 1698431365
transform 1 0 146384 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1037
timestamp 1698431365
transform 1 0 154224 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1038
timestamp 1698431365
transform 1 0 162064 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1039
timestamp 1698431365
transform 1 0 169904 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1040
timestamp 1698431365
transform 1 0 177744 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1041
timestamp 1698431365
transform 1 0 185584 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1042
timestamp 1698431365
transform 1 0 193424 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1043
timestamp 1698431365
transform 1 0 201264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1044
timestamp 1698431365
transform 1 0 209104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_1045
timestamp 1698431365
transform 1 0 216944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1046
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1047
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1048
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1049
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1050
timestamp 1698431365
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1051
timestamp 1698431365
transform 1 0 48384 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1052
timestamp 1698431365
transform 1 0 56224 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1053
timestamp 1698431365
transform 1 0 64064 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1054
timestamp 1698431365
transform 1 0 71904 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1055
timestamp 1698431365
transform 1 0 79744 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1056
timestamp 1698431365
transform 1 0 87584 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1057
timestamp 1698431365
transform 1 0 95424 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1058
timestamp 1698431365
transform 1 0 103264 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1059
timestamp 1698431365
transform 1 0 111104 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1060
timestamp 1698431365
transform 1 0 118944 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1061
timestamp 1698431365
transform 1 0 126784 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1062
timestamp 1698431365
transform 1 0 134624 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1063
timestamp 1698431365
transform 1 0 142464 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1064
timestamp 1698431365
transform 1 0 150304 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1065
timestamp 1698431365
transform 1 0 158144 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1066
timestamp 1698431365
transform 1 0 165984 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1067
timestamp 1698431365
transform 1 0 173824 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1068
timestamp 1698431365
transform 1 0 181664 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1069
timestamp 1698431365
transform 1 0 189504 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1070
timestamp 1698431365
transform 1 0 197344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1071
timestamp 1698431365
transform 1 0 205184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_1072
timestamp 1698431365
transform 1 0 213024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1073
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1074
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1075
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1076
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1077
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1078
timestamp 1698431365
transform 1 0 44464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1079
timestamp 1698431365
transform 1 0 52304 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1080
timestamp 1698431365
transform 1 0 60144 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1081
timestamp 1698431365
transform 1 0 67984 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1082
timestamp 1698431365
transform 1 0 75824 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1083
timestamp 1698431365
transform 1 0 83664 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1084
timestamp 1698431365
transform 1 0 91504 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1085
timestamp 1698431365
transform 1 0 99344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1086
timestamp 1698431365
transform 1 0 107184 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1087
timestamp 1698431365
transform 1 0 115024 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1088
timestamp 1698431365
transform 1 0 122864 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1089
timestamp 1698431365
transform 1 0 130704 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1090
timestamp 1698431365
transform 1 0 138544 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1091
timestamp 1698431365
transform 1 0 146384 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1092
timestamp 1698431365
transform 1 0 154224 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1093
timestamp 1698431365
transform 1 0 162064 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1094
timestamp 1698431365
transform 1 0 169904 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1095
timestamp 1698431365
transform 1 0 177744 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1096
timestamp 1698431365
transform 1 0 185584 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1097
timestamp 1698431365
transform 1 0 193424 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1098
timestamp 1698431365
transform 1 0 201264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1099
timestamp 1698431365
transform 1 0 209104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_1100
timestamp 1698431365
transform 1 0 216944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1101
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1102
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1103
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1104
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1105
timestamp 1698431365
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1106
timestamp 1698431365
transform 1 0 48384 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1107
timestamp 1698431365
transform 1 0 56224 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1108
timestamp 1698431365
transform 1 0 64064 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1109
timestamp 1698431365
transform 1 0 71904 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1110
timestamp 1698431365
transform 1 0 79744 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1111
timestamp 1698431365
transform 1 0 87584 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1112
timestamp 1698431365
transform 1 0 95424 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1113
timestamp 1698431365
transform 1 0 103264 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1114
timestamp 1698431365
transform 1 0 111104 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1115
timestamp 1698431365
transform 1 0 118944 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1116
timestamp 1698431365
transform 1 0 126784 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1117
timestamp 1698431365
transform 1 0 134624 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1118
timestamp 1698431365
transform 1 0 142464 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1119
timestamp 1698431365
transform 1 0 150304 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1120
timestamp 1698431365
transform 1 0 158144 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1121
timestamp 1698431365
transform 1 0 165984 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1122
timestamp 1698431365
transform 1 0 173824 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1123
timestamp 1698431365
transform 1 0 181664 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1124
timestamp 1698431365
transform 1 0 189504 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1125
timestamp 1698431365
transform 1 0 197344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1126
timestamp 1698431365
transform 1 0 205184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_1127
timestamp 1698431365
transform 1 0 213024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1128
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1129
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1130
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1131
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1132
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1133
timestamp 1698431365
transform 1 0 44464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1134
timestamp 1698431365
transform 1 0 52304 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1135
timestamp 1698431365
transform 1 0 60144 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1136
timestamp 1698431365
transform 1 0 67984 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1137
timestamp 1698431365
transform 1 0 75824 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1138
timestamp 1698431365
transform 1 0 83664 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1139
timestamp 1698431365
transform 1 0 91504 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1140
timestamp 1698431365
transform 1 0 99344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1141
timestamp 1698431365
transform 1 0 107184 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1142
timestamp 1698431365
transform 1 0 115024 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1143
timestamp 1698431365
transform 1 0 122864 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1144
timestamp 1698431365
transform 1 0 130704 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1145
timestamp 1698431365
transform 1 0 138544 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1146
timestamp 1698431365
transform 1 0 146384 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1147
timestamp 1698431365
transform 1 0 154224 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1148
timestamp 1698431365
transform 1 0 162064 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1149
timestamp 1698431365
transform 1 0 169904 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1150
timestamp 1698431365
transform 1 0 177744 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1151
timestamp 1698431365
transform 1 0 185584 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1152
timestamp 1698431365
transform 1 0 193424 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1153
timestamp 1698431365
transform 1 0 201264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1154
timestamp 1698431365
transform 1 0 209104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_1155
timestamp 1698431365
transform 1 0 216944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1156
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1157
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1158
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1159
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1160
timestamp 1698431365
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1161
timestamp 1698431365
transform 1 0 48384 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1162
timestamp 1698431365
transform 1 0 56224 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1163
timestamp 1698431365
transform 1 0 64064 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1164
timestamp 1698431365
transform 1 0 71904 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1165
timestamp 1698431365
transform 1 0 79744 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1166
timestamp 1698431365
transform 1 0 87584 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1167
timestamp 1698431365
transform 1 0 95424 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1168
timestamp 1698431365
transform 1 0 103264 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1169
timestamp 1698431365
transform 1 0 111104 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1170
timestamp 1698431365
transform 1 0 118944 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1171
timestamp 1698431365
transform 1 0 126784 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1172
timestamp 1698431365
transform 1 0 134624 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1173
timestamp 1698431365
transform 1 0 142464 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1174
timestamp 1698431365
transform 1 0 150304 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1175
timestamp 1698431365
transform 1 0 158144 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1176
timestamp 1698431365
transform 1 0 165984 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1177
timestamp 1698431365
transform 1 0 173824 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1178
timestamp 1698431365
transform 1 0 181664 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1179
timestamp 1698431365
transform 1 0 189504 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1180
timestamp 1698431365
transform 1 0 197344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1181
timestamp 1698431365
transform 1 0 205184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_1182
timestamp 1698431365
transform 1 0 213024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1183
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1184
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1185
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1186
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1187
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1188
timestamp 1698431365
transform 1 0 44464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1189
timestamp 1698431365
transform 1 0 52304 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1190
timestamp 1698431365
transform 1 0 60144 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1191
timestamp 1698431365
transform 1 0 67984 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1192
timestamp 1698431365
transform 1 0 75824 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1193
timestamp 1698431365
transform 1 0 83664 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1194
timestamp 1698431365
transform 1 0 91504 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1195
timestamp 1698431365
transform 1 0 99344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1196
timestamp 1698431365
transform 1 0 107184 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1197
timestamp 1698431365
transform 1 0 115024 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1198
timestamp 1698431365
transform 1 0 122864 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1199
timestamp 1698431365
transform 1 0 130704 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1200
timestamp 1698431365
transform 1 0 138544 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1201
timestamp 1698431365
transform 1 0 146384 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1202
timestamp 1698431365
transform 1 0 154224 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1203
timestamp 1698431365
transform 1 0 162064 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1204
timestamp 1698431365
transform 1 0 169904 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1205
timestamp 1698431365
transform 1 0 177744 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1206
timestamp 1698431365
transform 1 0 185584 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1207
timestamp 1698431365
transform 1 0 193424 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1208
timestamp 1698431365
transform 1 0 201264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1209
timestamp 1698431365
transform 1 0 209104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_1210
timestamp 1698431365
transform 1 0 216944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1211
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1212
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1213
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1214
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1215
timestamp 1698431365
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1216
timestamp 1698431365
transform 1 0 48384 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1217
timestamp 1698431365
transform 1 0 56224 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1218
timestamp 1698431365
transform 1 0 64064 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1219
timestamp 1698431365
transform 1 0 71904 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1220
timestamp 1698431365
transform 1 0 79744 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1221
timestamp 1698431365
transform 1 0 87584 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1222
timestamp 1698431365
transform 1 0 95424 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1223
timestamp 1698431365
transform 1 0 103264 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1224
timestamp 1698431365
transform 1 0 111104 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1225
timestamp 1698431365
transform 1 0 118944 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1226
timestamp 1698431365
transform 1 0 126784 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1227
timestamp 1698431365
transform 1 0 134624 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1228
timestamp 1698431365
transform 1 0 142464 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1229
timestamp 1698431365
transform 1 0 150304 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1230
timestamp 1698431365
transform 1 0 158144 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1231
timestamp 1698431365
transform 1 0 165984 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1232
timestamp 1698431365
transform 1 0 173824 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1233
timestamp 1698431365
transform 1 0 181664 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1234
timestamp 1698431365
transform 1 0 189504 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1235
timestamp 1698431365
transform 1 0 197344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1236
timestamp 1698431365
transform 1 0 205184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_1237
timestamp 1698431365
transform 1 0 213024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1238
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1239
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1240
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1241
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1242
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1243
timestamp 1698431365
transform 1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1244
timestamp 1698431365
transform 1 0 52304 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1245
timestamp 1698431365
transform 1 0 60144 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1246
timestamp 1698431365
transform 1 0 67984 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1247
timestamp 1698431365
transform 1 0 75824 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1248
timestamp 1698431365
transform 1 0 83664 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1249
timestamp 1698431365
transform 1 0 91504 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1250
timestamp 1698431365
transform 1 0 99344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1251
timestamp 1698431365
transform 1 0 107184 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1252
timestamp 1698431365
transform 1 0 115024 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1253
timestamp 1698431365
transform 1 0 122864 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1254
timestamp 1698431365
transform 1 0 130704 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1255
timestamp 1698431365
transform 1 0 138544 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1256
timestamp 1698431365
transform 1 0 146384 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1257
timestamp 1698431365
transform 1 0 154224 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1258
timestamp 1698431365
transform 1 0 162064 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1259
timestamp 1698431365
transform 1 0 169904 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1260
timestamp 1698431365
transform 1 0 177744 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1261
timestamp 1698431365
transform 1 0 185584 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1262
timestamp 1698431365
transform 1 0 193424 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1263
timestamp 1698431365
transform 1 0 201264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1264
timestamp 1698431365
transform 1 0 209104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_1265
timestamp 1698431365
transform 1 0 216944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1266
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1267
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1268
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1269
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1270
timestamp 1698431365
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1271
timestamp 1698431365
transform 1 0 48384 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1272
timestamp 1698431365
transform 1 0 56224 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1273
timestamp 1698431365
transform 1 0 64064 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1274
timestamp 1698431365
transform 1 0 71904 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1275
timestamp 1698431365
transform 1 0 79744 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1276
timestamp 1698431365
transform 1 0 87584 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1277
timestamp 1698431365
transform 1 0 95424 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1278
timestamp 1698431365
transform 1 0 103264 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1279
timestamp 1698431365
transform 1 0 111104 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1280
timestamp 1698431365
transform 1 0 118944 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1281
timestamp 1698431365
transform 1 0 126784 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1282
timestamp 1698431365
transform 1 0 134624 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1283
timestamp 1698431365
transform 1 0 142464 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1284
timestamp 1698431365
transform 1 0 150304 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1285
timestamp 1698431365
transform 1 0 158144 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1286
timestamp 1698431365
transform 1 0 165984 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1287
timestamp 1698431365
transform 1 0 173824 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1288
timestamp 1698431365
transform 1 0 181664 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1289
timestamp 1698431365
transform 1 0 189504 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1290
timestamp 1698431365
transform 1 0 197344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1291
timestamp 1698431365
transform 1 0 205184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_1292
timestamp 1698431365
transform 1 0 213024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1293
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1294
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1295
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1296
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1297
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1298
timestamp 1698431365
transform 1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1299
timestamp 1698431365
transform 1 0 52304 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1300
timestamp 1698431365
transform 1 0 60144 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1301
timestamp 1698431365
transform 1 0 67984 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1302
timestamp 1698431365
transform 1 0 75824 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1303
timestamp 1698431365
transform 1 0 83664 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1304
timestamp 1698431365
transform 1 0 91504 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1305
timestamp 1698431365
transform 1 0 99344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1306
timestamp 1698431365
transform 1 0 107184 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1307
timestamp 1698431365
transform 1 0 115024 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1308
timestamp 1698431365
transform 1 0 122864 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1309
timestamp 1698431365
transform 1 0 130704 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1310
timestamp 1698431365
transform 1 0 138544 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1311
timestamp 1698431365
transform 1 0 146384 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1312
timestamp 1698431365
transform 1 0 154224 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1313
timestamp 1698431365
transform 1 0 162064 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1314
timestamp 1698431365
transform 1 0 169904 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1315
timestamp 1698431365
transform 1 0 177744 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1316
timestamp 1698431365
transform 1 0 185584 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1317
timestamp 1698431365
transform 1 0 193424 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1318
timestamp 1698431365
transform 1 0 201264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1319
timestamp 1698431365
transform 1 0 209104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_1320
timestamp 1698431365
transform 1 0 216944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1321
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1322
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1323
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1324
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1325
timestamp 1698431365
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1326
timestamp 1698431365
transform 1 0 48384 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1327
timestamp 1698431365
transform 1 0 56224 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1328
timestamp 1698431365
transform 1 0 64064 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1329
timestamp 1698431365
transform 1 0 71904 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1330
timestamp 1698431365
transform 1 0 79744 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1331
timestamp 1698431365
transform 1 0 87584 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1332
timestamp 1698431365
transform 1 0 95424 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1333
timestamp 1698431365
transform 1 0 103264 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1334
timestamp 1698431365
transform 1 0 111104 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1335
timestamp 1698431365
transform 1 0 118944 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1336
timestamp 1698431365
transform 1 0 126784 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1337
timestamp 1698431365
transform 1 0 134624 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1338
timestamp 1698431365
transform 1 0 142464 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1339
timestamp 1698431365
transform 1 0 150304 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1340
timestamp 1698431365
transform 1 0 158144 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1341
timestamp 1698431365
transform 1 0 165984 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1342
timestamp 1698431365
transform 1 0 173824 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1343
timestamp 1698431365
transform 1 0 181664 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1344
timestamp 1698431365
transform 1 0 189504 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1345
timestamp 1698431365
transform 1 0 197344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1346
timestamp 1698431365
transform 1 0 205184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_1347
timestamp 1698431365
transform 1 0 213024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1348
timestamp 1698431365
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1349
timestamp 1698431365
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1350
timestamp 1698431365
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1351
timestamp 1698431365
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1352
timestamp 1698431365
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1353
timestamp 1698431365
transform 1 0 44464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1354
timestamp 1698431365
transform 1 0 52304 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1355
timestamp 1698431365
transform 1 0 60144 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1356
timestamp 1698431365
transform 1 0 67984 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1357
timestamp 1698431365
transform 1 0 75824 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1358
timestamp 1698431365
transform 1 0 83664 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1359
timestamp 1698431365
transform 1 0 91504 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1360
timestamp 1698431365
transform 1 0 99344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1361
timestamp 1698431365
transform 1 0 107184 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1362
timestamp 1698431365
transform 1 0 115024 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1363
timestamp 1698431365
transform 1 0 122864 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1364
timestamp 1698431365
transform 1 0 130704 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1365
timestamp 1698431365
transform 1 0 138544 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1366
timestamp 1698431365
transform 1 0 146384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1367
timestamp 1698431365
transform 1 0 154224 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1368
timestamp 1698431365
transform 1 0 162064 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1369
timestamp 1698431365
transform 1 0 169904 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1370
timestamp 1698431365
transform 1 0 177744 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1371
timestamp 1698431365
transform 1 0 185584 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1372
timestamp 1698431365
transform 1 0 193424 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1373
timestamp 1698431365
transform 1 0 201264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1374
timestamp 1698431365
transform 1 0 209104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_1375
timestamp 1698431365
transform 1 0 216944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1376
timestamp 1698431365
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1377
timestamp 1698431365
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1378
timestamp 1698431365
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1379
timestamp 1698431365
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1380
timestamp 1698431365
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1381
timestamp 1698431365
transform 1 0 48384 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1382
timestamp 1698431365
transform 1 0 56224 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1383
timestamp 1698431365
transform 1 0 64064 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1384
timestamp 1698431365
transform 1 0 71904 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1385
timestamp 1698431365
transform 1 0 79744 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1386
timestamp 1698431365
transform 1 0 87584 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1387
timestamp 1698431365
transform 1 0 95424 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1388
timestamp 1698431365
transform 1 0 103264 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1389
timestamp 1698431365
transform 1 0 111104 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1390
timestamp 1698431365
transform 1 0 118944 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1391
timestamp 1698431365
transform 1 0 126784 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1392
timestamp 1698431365
transform 1 0 134624 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1393
timestamp 1698431365
transform 1 0 142464 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1394
timestamp 1698431365
transform 1 0 150304 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1395
timestamp 1698431365
transform 1 0 158144 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1396
timestamp 1698431365
transform 1 0 165984 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1397
timestamp 1698431365
transform 1 0 173824 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1398
timestamp 1698431365
transform 1 0 181664 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1399
timestamp 1698431365
transform 1 0 189504 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1400
timestamp 1698431365
transform 1 0 197344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1401
timestamp 1698431365
transform 1 0 205184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_1402
timestamp 1698431365
transform 1 0 213024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1403
timestamp 1698431365
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1404
timestamp 1698431365
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1405
timestamp 1698431365
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1406
timestamp 1698431365
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1407
timestamp 1698431365
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1408
timestamp 1698431365
transform 1 0 44464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1409
timestamp 1698431365
transform 1 0 52304 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1410
timestamp 1698431365
transform 1 0 60144 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1411
timestamp 1698431365
transform 1 0 67984 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1412
timestamp 1698431365
transform 1 0 75824 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1413
timestamp 1698431365
transform 1 0 83664 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1414
timestamp 1698431365
transform 1 0 91504 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1415
timestamp 1698431365
transform 1 0 99344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1416
timestamp 1698431365
transform 1 0 107184 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1417
timestamp 1698431365
transform 1 0 115024 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1418
timestamp 1698431365
transform 1 0 122864 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1419
timestamp 1698431365
transform 1 0 130704 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1420
timestamp 1698431365
transform 1 0 138544 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1421
timestamp 1698431365
transform 1 0 146384 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1422
timestamp 1698431365
transform 1 0 154224 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1423
timestamp 1698431365
transform 1 0 162064 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1424
timestamp 1698431365
transform 1 0 169904 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1425
timestamp 1698431365
transform 1 0 177744 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1426
timestamp 1698431365
transform 1 0 185584 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1427
timestamp 1698431365
transform 1 0 193424 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1428
timestamp 1698431365
transform 1 0 201264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1429
timestamp 1698431365
transform 1 0 209104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_1430
timestamp 1698431365
transform 1 0 216944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1431
timestamp 1698431365
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1432
timestamp 1698431365
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1433
timestamp 1698431365
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1434
timestamp 1698431365
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1435
timestamp 1698431365
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1436
timestamp 1698431365
transform 1 0 48384 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1437
timestamp 1698431365
transform 1 0 56224 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1438
timestamp 1698431365
transform 1 0 64064 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1439
timestamp 1698431365
transform 1 0 71904 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1440
timestamp 1698431365
transform 1 0 79744 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1441
timestamp 1698431365
transform 1 0 87584 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1442
timestamp 1698431365
transform 1 0 95424 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1443
timestamp 1698431365
transform 1 0 103264 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1444
timestamp 1698431365
transform 1 0 111104 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1445
timestamp 1698431365
transform 1 0 118944 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1446
timestamp 1698431365
transform 1 0 126784 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1447
timestamp 1698431365
transform 1 0 134624 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1448
timestamp 1698431365
transform 1 0 142464 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1449
timestamp 1698431365
transform 1 0 150304 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1450
timestamp 1698431365
transform 1 0 158144 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1451
timestamp 1698431365
transform 1 0 165984 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1452
timestamp 1698431365
transform 1 0 173824 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1453
timestamp 1698431365
transform 1 0 181664 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1454
timestamp 1698431365
transform 1 0 189504 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1455
timestamp 1698431365
transform 1 0 197344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1456
timestamp 1698431365
transform 1 0 205184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_1457
timestamp 1698431365
transform 1 0 213024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1458
timestamp 1698431365
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1459
timestamp 1698431365
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1460
timestamp 1698431365
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1461
timestamp 1698431365
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1462
timestamp 1698431365
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1463
timestamp 1698431365
transform 1 0 44464 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1464
timestamp 1698431365
transform 1 0 52304 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1465
timestamp 1698431365
transform 1 0 60144 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1466
timestamp 1698431365
transform 1 0 67984 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1467
timestamp 1698431365
transform 1 0 75824 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1468
timestamp 1698431365
transform 1 0 83664 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1469
timestamp 1698431365
transform 1 0 91504 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1470
timestamp 1698431365
transform 1 0 99344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1471
timestamp 1698431365
transform 1 0 107184 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1472
timestamp 1698431365
transform 1 0 115024 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1473
timestamp 1698431365
transform 1 0 122864 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1474
timestamp 1698431365
transform 1 0 130704 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1475
timestamp 1698431365
transform 1 0 138544 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1476
timestamp 1698431365
transform 1 0 146384 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1477
timestamp 1698431365
transform 1 0 154224 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1478
timestamp 1698431365
transform 1 0 162064 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1479
timestamp 1698431365
transform 1 0 169904 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1480
timestamp 1698431365
transform 1 0 177744 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1481
timestamp 1698431365
transform 1 0 185584 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1482
timestamp 1698431365
transform 1 0 193424 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1483
timestamp 1698431365
transform 1 0 201264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1484
timestamp 1698431365
transform 1 0 209104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_1485
timestamp 1698431365
transform 1 0 216944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1486
timestamp 1698431365
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1487
timestamp 1698431365
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1488
timestamp 1698431365
transform 1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1489
timestamp 1698431365
transform 1 0 32704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1490
timestamp 1698431365
transform 1 0 40544 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1491
timestamp 1698431365
transform 1 0 48384 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1492
timestamp 1698431365
transform 1 0 56224 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1493
timestamp 1698431365
transform 1 0 64064 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1494
timestamp 1698431365
transform 1 0 71904 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1495
timestamp 1698431365
transform 1 0 79744 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1496
timestamp 1698431365
transform 1 0 87584 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1497
timestamp 1698431365
transform 1 0 95424 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1498
timestamp 1698431365
transform 1 0 103264 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1499
timestamp 1698431365
transform 1 0 111104 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1500
timestamp 1698431365
transform 1 0 118944 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1501
timestamp 1698431365
transform 1 0 126784 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1502
timestamp 1698431365
transform 1 0 134624 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1503
timestamp 1698431365
transform 1 0 142464 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1504
timestamp 1698431365
transform 1 0 150304 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1505
timestamp 1698431365
transform 1 0 158144 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1506
timestamp 1698431365
transform 1 0 165984 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1507
timestamp 1698431365
transform 1 0 173824 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1508
timestamp 1698431365
transform 1 0 181664 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1509
timestamp 1698431365
transform 1 0 189504 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1510
timestamp 1698431365
transform 1 0 197344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1511
timestamp 1698431365
transform 1 0 205184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_1512
timestamp 1698431365
transform 1 0 213024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1513
timestamp 1698431365
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1514
timestamp 1698431365
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1515
timestamp 1698431365
transform 1 0 20944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1516
timestamp 1698431365
transform 1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1517
timestamp 1698431365
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1518
timestamp 1698431365
transform 1 0 44464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1519
timestamp 1698431365
transform 1 0 52304 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1520
timestamp 1698431365
transform 1 0 60144 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1521
timestamp 1698431365
transform 1 0 67984 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1522
timestamp 1698431365
transform 1 0 75824 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1523
timestamp 1698431365
transform 1 0 83664 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1524
timestamp 1698431365
transform 1 0 91504 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1525
timestamp 1698431365
transform 1 0 99344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1526
timestamp 1698431365
transform 1 0 107184 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1527
timestamp 1698431365
transform 1 0 115024 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1528
timestamp 1698431365
transform 1 0 122864 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1529
timestamp 1698431365
transform 1 0 130704 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1530
timestamp 1698431365
transform 1 0 138544 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1531
timestamp 1698431365
transform 1 0 146384 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1532
timestamp 1698431365
transform 1 0 154224 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1533
timestamp 1698431365
transform 1 0 162064 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1534
timestamp 1698431365
transform 1 0 169904 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1535
timestamp 1698431365
transform 1 0 177744 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1536
timestamp 1698431365
transform 1 0 185584 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1537
timestamp 1698431365
transform 1 0 193424 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1538
timestamp 1698431365
transform 1 0 201264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1539
timestamp 1698431365
transform 1 0 209104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_1540
timestamp 1698431365
transform 1 0 216944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1541
timestamp 1698431365
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1542
timestamp 1698431365
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1543
timestamp 1698431365
transform 1 0 24864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1544
timestamp 1698431365
transform 1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1545
timestamp 1698431365
transform 1 0 40544 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1546
timestamp 1698431365
transform 1 0 48384 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1547
timestamp 1698431365
transform 1 0 56224 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1548
timestamp 1698431365
transform 1 0 64064 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1549
timestamp 1698431365
transform 1 0 71904 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1550
timestamp 1698431365
transform 1 0 79744 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1551
timestamp 1698431365
transform 1 0 87584 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1552
timestamp 1698431365
transform 1 0 95424 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1553
timestamp 1698431365
transform 1 0 103264 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1554
timestamp 1698431365
transform 1 0 111104 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1555
timestamp 1698431365
transform 1 0 118944 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1556
timestamp 1698431365
transform 1 0 126784 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1557
timestamp 1698431365
transform 1 0 134624 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1558
timestamp 1698431365
transform 1 0 142464 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1559
timestamp 1698431365
transform 1 0 150304 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1560
timestamp 1698431365
transform 1 0 158144 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1561
timestamp 1698431365
transform 1 0 165984 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1562
timestamp 1698431365
transform 1 0 173824 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1563
timestamp 1698431365
transform 1 0 181664 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1564
timestamp 1698431365
transform 1 0 189504 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1565
timestamp 1698431365
transform 1 0 197344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1566
timestamp 1698431365
transform 1 0 205184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_1567
timestamp 1698431365
transform 1 0 213024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1568
timestamp 1698431365
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1569
timestamp 1698431365
transform 1 0 13104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1570
timestamp 1698431365
transform 1 0 20944 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1571
timestamp 1698431365
transform 1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1572
timestamp 1698431365
transform 1 0 36624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1573
timestamp 1698431365
transform 1 0 44464 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1574
timestamp 1698431365
transform 1 0 52304 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1575
timestamp 1698431365
transform 1 0 60144 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1576
timestamp 1698431365
transform 1 0 67984 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1577
timestamp 1698431365
transform 1 0 75824 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1578
timestamp 1698431365
transform 1 0 83664 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1579
timestamp 1698431365
transform 1 0 91504 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1580
timestamp 1698431365
transform 1 0 99344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1581
timestamp 1698431365
transform 1 0 107184 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1582
timestamp 1698431365
transform 1 0 115024 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1583
timestamp 1698431365
transform 1 0 122864 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1584
timestamp 1698431365
transform 1 0 130704 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1585
timestamp 1698431365
transform 1 0 138544 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1586
timestamp 1698431365
transform 1 0 146384 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1587
timestamp 1698431365
transform 1 0 154224 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1588
timestamp 1698431365
transform 1 0 162064 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1589
timestamp 1698431365
transform 1 0 169904 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1590
timestamp 1698431365
transform 1 0 177744 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1591
timestamp 1698431365
transform 1 0 185584 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1592
timestamp 1698431365
transform 1 0 193424 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1593
timestamp 1698431365
transform 1 0 201264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1594
timestamp 1698431365
transform 1 0 209104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_1595
timestamp 1698431365
transform 1 0 216944 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1596
timestamp 1698431365
transform 1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1597
timestamp 1698431365
transform 1 0 17024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1598
timestamp 1698431365
transform 1 0 24864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1599
timestamp 1698431365
transform 1 0 32704 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1600
timestamp 1698431365
transform 1 0 40544 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1601
timestamp 1698431365
transform 1 0 48384 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1602
timestamp 1698431365
transform 1 0 56224 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1603
timestamp 1698431365
transform 1 0 64064 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1604
timestamp 1698431365
transform 1 0 71904 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1605
timestamp 1698431365
transform 1 0 79744 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1606
timestamp 1698431365
transform 1 0 87584 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1607
timestamp 1698431365
transform 1 0 95424 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1608
timestamp 1698431365
transform 1 0 103264 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1609
timestamp 1698431365
transform 1 0 111104 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1610
timestamp 1698431365
transform 1 0 118944 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1611
timestamp 1698431365
transform 1 0 126784 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1612
timestamp 1698431365
transform 1 0 134624 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1613
timestamp 1698431365
transform 1 0 142464 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1614
timestamp 1698431365
transform 1 0 150304 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1615
timestamp 1698431365
transform 1 0 158144 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1616
timestamp 1698431365
transform 1 0 165984 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1617
timestamp 1698431365
transform 1 0 173824 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1618
timestamp 1698431365
transform 1 0 181664 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1619
timestamp 1698431365
transform 1 0 189504 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1620
timestamp 1698431365
transform 1 0 197344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1621
timestamp 1698431365
transform 1 0 205184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_1622
timestamp 1698431365
transform 1 0 213024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1623
timestamp 1698431365
transform 1 0 5152 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1624
timestamp 1698431365
transform 1 0 8960 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1625
timestamp 1698431365
transform 1 0 12768 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1626
timestamp 1698431365
transform 1 0 16576 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1627
timestamp 1698431365
transform 1 0 20384 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1628
timestamp 1698431365
transform 1 0 24192 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1629
timestamp 1698431365
transform 1 0 28000 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1630
timestamp 1698431365
transform 1 0 31808 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1631
timestamp 1698431365
transform 1 0 35616 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1632
timestamp 1698431365
transform 1 0 39424 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1633
timestamp 1698431365
transform 1 0 43232 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1634
timestamp 1698431365
transform 1 0 47040 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1635
timestamp 1698431365
transform 1 0 50848 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1636
timestamp 1698431365
transform 1 0 54656 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1637
timestamp 1698431365
transform 1 0 58464 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1638
timestamp 1698431365
transform 1 0 62272 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1639
timestamp 1698431365
transform 1 0 66080 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1640
timestamp 1698431365
transform 1 0 69888 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1641
timestamp 1698431365
transform 1 0 73696 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1642
timestamp 1698431365
transform 1 0 77504 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1643
timestamp 1698431365
transform 1 0 81312 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1644
timestamp 1698431365
transform 1 0 85120 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1645
timestamp 1698431365
transform 1 0 88928 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1646
timestamp 1698431365
transform 1 0 92736 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1647
timestamp 1698431365
transform 1 0 96544 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1648
timestamp 1698431365
transform 1 0 100352 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1649
timestamp 1698431365
transform 1 0 104160 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1650
timestamp 1698431365
transform 1 0 107968 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1651
timestamp 1698431365
transform 1 0 111776 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1652
timestamp 1698431365
transform 1 0 115584 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1653
timestamp 1698431365
transform 1 0 119392 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1654
timestamp 1698431365
transform 1 0 123200 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1655
timestamp 1698431365
transform 1 0 127008 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1656
timestamp 1698431365
transform 1 0 130816 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1657
timestamp 1698431365
transform 1 0 134624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1658
timestamp 1698431365
transform 1 0 138432 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1659
timestamp 1698431365
transform 1 0 142240 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1660
timestamp 1698431365
transform 1 0 146048 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1661
timestamp 1698431365
transform 1 0 149856 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1662
timestamp 1698431365
transform 1 0 153664 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1663
timestamp 1698431365
transform 1 0 157472 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1664
timestamp 1698431365
transform 1 0 161280 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1665
timestamp 1698431365
transform 1 0 165088 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1666
timestamp 1698431365
transform 1 0 168896 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1667
timestamp 1698431365
transform 1 0 172704 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1668
timestamp 1698431365
transform 1 0 176512 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1669
timestamp 1698431365
transform 1 0 180320 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1670
timestamp 1698431365
transform 1 0 184128 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1671
timestamp 1698431365
transform 1 0 187936 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1672
timestamp 1698431365
transform 1 0 191744 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1673
timestamp 1698431365
transform 1 0 195552 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1674
timestamp 1698431365
transform 1 0 199360 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1675
timestamp 1698431365
transform 1 0 203168 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1676
timestamp 1698431365
transform 1 0 206976 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1677
timestamp 1698431365
transform 1 0 210784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_1678
timestamp 1698431365
transform 1 0 214592 0 1 45472
box -86 -86 310 870
<< labels >>
flabel metal2 s 27776 0 27888 800 0 FreeSans 448 90 0 0 A_all[0]
port 0 nsew signal tristate
flabel metal2 s 30464 0 30576 800 0 FreeSans 448 90 0 0 A_all[1]
port 1 nsew signal tristate
flabel metal2 s 33152 0 33264 800 0 FreeSans 448 90 0 0 A_all[2]
port 2 nsew signal tristate
flabel metal2 s 35840 0 35952 800 0 FreeSans 448 90 0 0 A_all[3]
port 3 nsew signal tristate
flabel metal2 s 38528 0 38640 800 0 FreeSans 448 90 0 0 A_all[4]
port 4 nsew signal tristate
flabel metal2 s 41216 0 41328 800 0 FreeSans 448 90 0 0 A_all[5]
port 5 nsew signal tristate
flabel metal2 s 43904 0 44016 800 0 FreeSans 448 90 0 0 A_all[6]
port 6 nsew signal tristate
flabel metal2 s 46592 0 46704 800 0 FreeSans 448 90 0 0 A_all[7]
port 7 nsew signal tristate
flabel metal2 s 49280 0 49392 800 0 FreeSans 448 90 0 0 A_all[8]
port 8 nsew signal tristate
flabel metal2 s 3584 0 3696 800 0 FreeSans 448 90 0 0 CEN_all
port 9 nsew signal tristate
flabel metal2 s 51968 0 52080 800 0 FreeSans 448 90 0 0 D_all[0]
port 10 nsew signal tristate
flabel metal2 s 54656 0 54768 800 0 FreeSans 448 90 0 0 D_all[1]
port 11 nsew signal tristate
flabel metal2 s 57344 0 57456 800 0 FreeSans 448 90 0 0 D_all[2]
port 12 nsew signal tristate
flabel metal2 s 60032 0 60144 800 0 FreeSans 448 90 0 0 D_all[3]
port 13 nsew signal tristate
flabel metal2 s 62720 0 62832 800 0 FreeSans 448 90 0 0 D_all[4]
port 14 nsew signal tristate
flabel metal2 s 65408 0 65520 800 0 FreeSans 448 90 0 0 D_all[5]
port 15 nsew signal tristate
flabel metal2 s 68096 0 68208 800 0 FreeSans 448 90 0 0 D_all[6]
port 16 nsew signal tristate
flabel metal2 s 70784 0 70896 800 0 FreeSans 448 90 0 0 D_all[7]
port 17 nsew signal tristate
flabel metal2 s 73472 0 73584 800 0 FreeSans 448 90 0 0 GWEN_0
port 18 nsew signal tristate
flabel metal2 s 76160 0 76272 800 0 FreeSans 448 90 0 0 GWEN_1
port 19 nsew signal tristate
flabel metal2 s 78848 0 78960 800 0 FreeSans 448 90 0 0 GWEN_2
port 20 nsew signal tristate
flabel metal2 s 81536 0 81648 800 0 FreeSans 448 90 0 0 GWEN_3
port 21 nsew signal tristate
flabel metal2 s 84224 0 84336 800 0 FreeSans 448 90 0 0 GWEN_4
port 22 nsew signal tristate
flabel metal2 s 86912 0 87024 800 0 FreeSans 448 90 0 0 GWEN_5
port 23 nsew signal tristate
flabel metal2 s 148064 49200 148176 50000 0 FreeSans 448 90 0 0 GWEN_6
port 24 nsew signal tristate
flabel metal2 s 152096 49200 152208 50000 0 FreeSans 448 90 0 0 GWEN_7
port 25 nsew signal tristate
flabel metal2 s 89600 0 89712 800 0 FreeSans 448 90 0 0 Q0[0]
port 26 nsew signal input
flabel metal2 s 92288 0 92400 800 0 FreeSans 448 90 0 0 Q0[1]
port 27 nsew signal input
flabel metal2 s 94976 0 95088 800 0 FreeSans 448 90 0 0 Q0[2]
port 28 nsew signal input
flabel metal2 s 97664 0 97776 800 0 FreeSans 448 90 0 0 Q0[3]
port 29 nsew signal input
flabel metal2 s 100352 0 100464 800 0 FreeSans 448 90 0 0 Q0[4]
port 30 nsew signal input
flabel metal2 s 103040 0 103152 800 0 FreeSans 448 90 0 0 Q0[5]
port 31 nsew signal input
flabel metal2 s 105728 0 105840 800 0 FreeSans 448 90 0 0 Q0[6]
port 32 nsew signal input
flabel metal2 s 108416 0 108528 800 0 FreeSans 448 90 0 0 Q0[7]
port 33 nsew signal input
flabel metal2 s 111104 0 111216 800 0 FreeSans 448 90 0 0 Q1[0]
port 34 nsew signal input
flabel metal2 s 113792 0 113904 800 0 FreeSans 448 90 0 0 Q1[1]
port 35 nsew signal input
flabel metal2 s 116480 0 116592 800 0 FreeSans 448 90 0 0 Q1[2]
port 36 nsew signal input
flabel metal2 s 119168 0 119280 800 0 FreeSans 448 90 0 0 Q1[3]
port 37 nsew signal input
flabel metal2 s 121856 0 121968 800 0 FreeSans 448 90 0 0 Q1[4]
port 38 nsew signal input
flabel metal2 s 124544 0 124656 800 0 FreeSans 448 90 0 0 Q1[5]
port 39 nsew signal input
flabel metal2 s 127232 0 127344 800 0 FreeSans 448 90 0 0 Q1[6]
port 40 nsew signal input
flabel metal2 s 129920 0 130032 800 0 FreeSans 448 90 0 0 Q1[7]
port 41 nsew signal input
flabel metal2 s 132608 0 132720 800 0 FreeSans 448 90 0 0 Q2[0]
port 42 nsew signal input
flabel metal2 s 135296 0 135408 800 0 FreeSans 448 90 0 0 Q2[1]
port 43 nsew signal input
flabel metal2 s 137984 0 138096 800 0 FreeSans 448 90 0 0 Q2[2]
port 44 nsew signal input
flabel metal2 s 140672 0 140784 800 0 FreeSans 448 90 0 0 Q2[3]
port 45 nsew signal input
flabel metal2 s 143360 0 143472 800 0 FreeSans 448 90 0 0 Q2[4]
port 46 nsew signal input
flabel metal2 s 146048 0 146160 800 0 FreeSans 448 90 0 0 Q2[5]
port 47 nsew signal input
flabel metal2 s 148736 0 148848 800 0 FreeSans 448 90 0 0 Q2[6]
port 48 nsew signal input
flabel metal2 s 151424 0 151536 800 0 FreeSans 448 90 0 0 Q2[7]
port 49 nsew signal input
flabel metal2 s 154112 0 154224 800 0 FreeSans 448 90 0 0 Q3[0]
port 50 nsew signal input
flabel metal2 s 156800 0 156912 800 0 FreeSans 448 90 0 0 Q3[1]
port 51 nsew signal input
flabel metal2 s 159488 0 159600 800 0 FreeSans 448 90 0 0 Q3[2]
port 52 nsew signal input
flabel metal2 s 162176 0 162288 800 0 FreeSans 448 90 0 0 Q3[3]
port 53 nsew signal input
flabel metal2 s 164864 0 164976 800 0 FreeSans 448 90 0 0 Q3[4]
port 54 nsew signal input
flabel metal2 s 167552 0 167664 800 0 FreeSans 448 90 0 0 Q3[5]
port 55 nsew signal input
flabel metal2 s 170240 0 170352 800 0 FreeSans 448 90 0 0 Q3[6]
port 56 nsew signal input
flabel metal2 s 172928 0 173040 800 0 FreeSans 448 90 0 0 Q3[7]
port 57 nsew signal input
flabel metal2 s 175616 0 175728 800 0 FreeSans 448 90 0 0 Q4[0]
port 58 nsew signal input
flabel metal2 s 178304 0 178416 800 0 FreeSans 448 90 0 0 Q4[1]
port 59 nsew signal input
flabel metal2 s 180992 0 181104 800 0 FreeSans 448 90 0 0 Q4[2]
port 60 nsew signal input
flabel metal2 s 183680 0 183792 800 0 FreeSans 448 90 0 0 Q4[3]
port 61 nsew signal input
flabel metal2 s 186368 0 186480 800 0 FreeSans 448 90 0 0 Q4[4]
port 62 nsew signal input
flabel metal2 s 189056 0 189168 800 0 FreeSans 448 90 0 0 Q4[5]
port 63 nsew signal input
flabel metal2 s 191744 0 191856 800 0 FreeSans 448 90 0 0 Q4[6]
port 64 nsew signal input
flabel metal2 s 194432 0 194544 800 0 FreeSans 448 90 0 0 Q4[7]
port 65 nsew signal input
flabel metal2 s 197120 0 197232 800 0 FreeSans 448 90 0 0 Q5[0]
port 66 nsew signal input
flabel metal2 s 199808 0 199920 800 0 FreeSans 448 90 0 0 Q5[1]
port 67 nsew signal input
flabel metal2 s 202496 0 202608 800 0 FreeSans 448 90 0 0 Q5[2]
port 68 nsew signal input
flabel metal2 s 205184 0 205296 800 0 FreeSans 448 90 0 0 Q5[3]
port 69 nsew signal input
flabel metal2 s 207872 0 207984 800 0 FreeSans 448 90 0 0 Q5[4]
port 70 nsew signal input
flabel metal2 s 210560 0 210672 800 0 FreeSans 448 90 0 0 Q5[5]
port 71 nsew signal input
flabel metal2 s 213248 0 213360 800 0 FreeSans 448 90 0 0 Q5[6]
port 72 nsew signal input
flabel metal2 s 215936 0 216048 800 0 FreeSans 448 90 0 0 Q5[7]
port 73 nsew signal input
flabel metal2 s 156128 49200 156240 50000 0 FreeSans 448 90 0 0 Q6[0]
port 74 nsew signal input
flabel metal2 s 160160 49200 160272 50000 0 FreeSans 448 90 0 0 Q6[1]
port 75 nsew signal input
flabel metal2 s 164192 49200 164304 50000 0 FreeSans 448 90 0 0 Q6[2]
port 76 nsew signal input
flabel metal2 s 168224 49200 168336 50000 0 FreeSans 448 90 0 0 Q6[3]
port 77 nsew signal input
flabel metal2 s 172256 49200 172368 50000 0 FreeSans 448 90 0 0 Q6[4]
port 78 nsew signal input
flabel metal2 s 176288 49200 176400 50000 0 FreeSans 448 90 0 0 Q6[5]
port 79 nsew signal input
flabel metal2 s 180320 49200 180432 50000 0 FreeSans 448 90 0 0 Q6[6]
port 80 nsew signal input
flabel metal2 s 184352 49200 184464 50000 0 FreeSans 448 90 0 0 Q6[7]
port 81 nsew signal input
flabel metal2 s 188384 49200 188496 50000 0 FreeSans 448 90 0 0 Q7[0]
port 82 nsew signal input
flabel metal2 s 192416 49200 192528 50000 0 FreeSans 448 90 0 0 Q7[1]
port 83 nsew signal input
flabel metal2 s 196448 49200 196560 50000 0 FreeSans 448 90 0 0 Q7[2]
port 84 nsew signal input
flabel metal2 s 200480 49200 200592 50000 0 FreeSans 448 90 0 0 Q7[3]
port 85 nsew signal input
flabel metal2 s 204512 49200 204624 50000 0 FreeSans 448 90 0 0 Q7[4]
port 86 nsew signal input
flabel metal2 s 208544 49200 208656 50000 0 FreeSans 448 90 0 0 Q7[5]
port 87 nsew signal input
flabel metal2 s 212576 49200 212688 50000 0 FreeSans 448 90 0 0 Q7[6]
port 88 nsew signal input
flabel metal2 s 216608 49200 216720 50000 0 FreeSans 448 90 0 0 Q7[7]
port 89 nsew signal input
flabel metal2 s 6272 0 6384 800 0 FreeSans 448 90 0 0 WEN_all[0]
port 90 nsew signal tristate
flabel metal2 s 8960 0 9072 800 0 FreeSans 448 90 0 0 WEN_all[1]
port 91 nsew signal tristate
flabel metal2 s 11648 0 11760 800 0 FreeSans 448 90 0 0 WEN_all[2]
port 92 nsew signal tristate
flabel metal2 s 14336 0 14448 800 0 FreeSans 448 90 0 0 WEN_all[3]
port 93 nsew signal tristate
flabel metal2 s 17024 0 17136 800 0 FreeSans 448 90 0 0 WEN_all[4]
port 94 nsew signal tristate
flabel metal2 s 19712 0 19824 800 0 FreeSans 448 90 0 0 WEN_all[5]
port 95 nsew signal tristate
flabel metal2 s 22400 0 22512 800 0 FreeSans 448 90 0 0 WEN_all[6]
port 96 nsew signal tristate
flabel metal2 s 25088 0 25200 800 0 FreeSans 448 90 0 0 WEN_all[7]
port 97 nsew signal tristate
flabel metal2 s 10976 49200 11088 50000 0 FreeSans 448 90 0 0 WEb_ram
port 98 nsew signal input
flabel metal2 s 15008 49200 15120 50000 0 FreeSans 448 90 0 0 bus_in[0]
port 99 nsew signal input
flabel metal2 s 19040 49200 19152 50000 0 FreeSans 448 90 0 0 bus_in[1]
port 100 nsew signal input
flabel metal2 s 23072 49200 23184 50000 0 FreeSans 448 90 0 0 bus_in[2]
port 101 nsew signal input
flabel metal2 s 27104 49200 27216 50000 0 FreeSans 448 90 0 0 bus_in[3]
port 102 nsew signal input
flabel metal2 s 31136 49200 31248 50000 0 FreeSans 448 90 0 0 bus_in[4]
port 103 nsew signal input
flabel metal2 s 35168 49200 35280 50000 0 FreeSans 448 90 0 0 bus_in[5]
port 104 nsew signal input
flabel metal2 s 39200 49200 39312 50000 0 FreeSans 448 90 0 0 bus_in[6]
port 105 nsew signal input
flabel metal2 s 43232 49200 43344 50000 0 FreeSans 448 90 0 0 bus_in[7]
port 106 nsew signal input
flabel metal2 s 47264 49200 47376 50000 0 FreeSans 448 90 0 0 bus_out[0]
port 107 nsew signal tristate
flabel metal2 s 51296 49200 51408 50000 0 FreeSans 448 90 0 0 bus_out[1]
port 108 nsew signal tristate
flabel metal2 s 55328 49200 55440 50000 0 FreeSans 448 90 0 0 bus_out[2]
port 109 nsew signal tristate
flabel metal2 s 59360 49200 59472 50000 0 FreeSans 448 90 0 0 bus_out[3]
port 110 nsew signal tristate
flabel metal2 s 63392 49200 63504 50000 0 FreeSans 448 90 0 0 bus_out[4]
port 111 nsew signal tristate
flabel metal2 s 67424 49200 67536 50000 0 FreeSans 448 90 0 0 bus_out[5]
port 112 nsew signal tristate
flabel metal2 s 71456 49200 71568 50000 0 FreeSans 448 90 0 0 bus_out[6]
port 113 nsew signal tristate
flabel metal2 s 75488 49200 75600 50000 0 FreeSans 448 90 0 0 bus_out[7]
port 114 nsew signal tristate
flabel metal2 s 79520 49200 79632 50000 0 FreeSans 448 90 0 0 ram_enabled
port 115 nsew signal input
flabel metal2 s 83552 49200 83664 50000 0 FreeSans 448 90 0 0 requested_addr[0]
port 116 nsew signal input
flabel metal2 s 123872 49200 123984 50000 0 FreeSans 448 90 0 0 requested_addr[10]
port 117 nsew signal input
flabel metal2 s 127904 49200 128016 50000 0 FreeSans 448 90 0 0 requested_addr[11]
port 118 nsew signal input
flabel metal2 s 131936 49200 132048 50000 0 FreeSans 448 90 0 0 requested_addr[12]
port 119 nsew signal input
flabel metal2 s 135968 49200 136080 50000 0 FreeSans 448 90 0 0 requested_addr[13]
port 120 nsew signal input
flabel metal2 s 140000 49200 140112 50000 0 FreeSans 448 90 0 0 requested_addr[14]
port 121 nsew signal input
flabel metal2 s 144032 49200 144144 50000 0 FreeSans 448 90 0 0 requested_addr[15]
port 122 nsew signal input
flabel metal2 s 87584 49200 87696 50000 0 FreeSans 448 90 0 0 requested_addr[1]
port 123 nsew signal input
flabel metal2 s 91616 49200 91728 50000 0 FreeSans 448 90 0 0 requested_addr[2]
port 124 nsew signal input
flabel metal2 s 95648 49200 95760 50000 0 FreeSans 448 90 0 0 requested_addr[3]
port 125 nsew signal input
flabel metal2 s 99680 49200 99792 50000 0 FreeSans 448 90 0 0 requested_addr[4]
port 126 nsew signal input
flabel metal2 s 103712 49200 103824 50000 0 FreeSans 448 90 0 0 requested_addr[5]
port 127 nsew signal input
flabel metal2 s 107744 49200 107856 50000 0 FreeSans 448 90 0 0 requested_addr[6]
port 128 nsew signal input
flabel metal2 s 111776 49200 111888 50000 0 FreeSans 448 90 0 0 requested_addr[7]
port 129 nsew signal input
flabel metal2 s 115808 49200 115920 50000 0 FreeSans 448 90 0 0 requested_addr[8]
port 130 nsew signal input
flabel metal2 s 119840 49200 119952 50000 0 FreeSans 448 90 0 0 requested_addr[9]
port 131 nsew signal input
flabel metal2 s 6944 49200 7056 50000 0 FreeSans 448 90 0 0 rst
port 132 nsew signal input
flabel metal4 s 4448 3076 4768 46316 0 FreeSans 1280 90 0 0 vdd
port 133 nsew power bidirectional
flabel metal4 s 35168 3076 35488 46316 0 FreeSans 1280 90 0 0 vdd
port 133 nsew power bidirectional
flabel metal4 s 65888 3076 66208 46316 0 FreeSans 1280 90 0 0 vdd
port 133 nsew power bidirectional
flabel metal4 s 96608 3076 96928 46316 0 FreeSans 1280 90 0 0 vdd
port 133 nsew power bidirectional
flabel metal4 s 127328 3076 127648 46316 0 FreeSans 1280 90 0 0 vdd
port 133 nsew power bidirectional
flabel metal4 s 158048 3076 158368 46316 0 FreeSans 1280 90 0 0 vdd
port 133 nsew power bidirectional
flabel metal4 s 188768 3076 189088 46316 0 FreeSans 1280 90 0 0 vdd
port 133 nsew power bidirectional
flabel metal4 s 19808 3076 20128 46316 0 FreeSans 1280 90 0 0 vss
port 134 nsew ground bidirectional
flabel metal4 s 50528 3076 50848 46316 0 FreeSans 1280 90 0 0 vss
port 134 nsew ground bidirectional
flabel metal4 s 81248 3076 81568 46316 0 FreeSans 1280 90 0 0 vss
port 134 nsew ground bidirectional
flabel metal4 s 111968 3076 112288 46316 0 FreeSans 1280 90 0 0 vss
port 134 nsew ground bidirectional
flabel metal4 s 142688 3076 143008 46316 0 FreeSans 1280 90 0 0 vss
port 134 nsew ground bidirectional
flabel metal4 s 173408 3076 173728 46316 0 FreeSans 1280 90 0 0 vss
port 134 nsew ground bidirectional
flabel metal4 s 204128 3076 204448 46316 0 FreeSans 1280 90 0 0 vss
port 134 nsew ground bidirectional
flabel metal2 s 2912 49200 3024 50000 0 FreeSans 448 90 0 0 wb_clk_i
port 135 nsew signal input
rlabel metal1 109984 46256 109984 46256 0 vdd
rlabel metal1 109984 45472 109984 45472 0 vss
rlabel metal2 27832 2198 27832 2198 0 A_all[0]
rlabel metal2 30520 1414 30520 1414 0 A_all[1]
rlabel metal2 33208 2198 33208 2198 0 A_all[2]
rlabel metal2 35896 2198 35896 2198 0 A_all[3]
rlabel metal2 38584 2086 38584 2086 0 A_all[4]
rlabel metal2 41272 2422 41272 2422 0 A_all[5]
rlabel metal2 43960 2198 43960 2198 0 A_all[6]
rlabel metal2 46648 2086 46648 2086 0 A_all[7]
rlabel metal2 49336 2422 49336 2422 0 A_all[8]
rlabel metal2 3640 2422 3640 2422 0 CEN_all
rlabel metal2 52024 2086 52024 2086 0 D_all[0]
rlabel metal2 54712 2086 54712 2086 0 D_all[1]
rlabel metal2 57400 2422 57400 2422 0 D_all[2]
rlabel metal2 60088 2198 60088 2198 0 D_all[3]
rlabel metal2 62776 2198 62776 2198 0 D_all[4]
rlabel metal3 67480 3528 67480 3528 0 D_all[5]
rlabel metal2 68152 2422 68152 2422 0 D_all[6]
rlabel metal2 70840 2086 70840 2086 0 D_all[7]
rlabel metal2 73528 2198 73528 2198 0 GWEN_0
rlabel metal2 76216 2422 76216 2422 0 GWEN_1
rlabel metal2 78904 2198 78904 2198 0 GWEN_2
rlabel metal2 81592 854 81592 854 0 GWEN_3
rlabel metal2 84280 2422 84280 2422 0 GWEN_4
rlabel metal2 86968 2086 86968 2086 0 GWEN_5
rlabel metal2 148120 47698 148120 47698 0 GWEN_6
rlabel metal2 152152 47306 152152 47306 0 GWEN_7
rlabel metal2 89656 2086 89656 2086 0 Q0[0]
rlabel metal2 92512 3416 92512 3416 0 Q0[1]
rlabel metal2 95032 2086 95032 2086 0 Q0[2]
rlabel metal2 97720 2086 97720 2086 0 Q0[3]
rlabel metal2 100352 3416 100352 3416 0 Q0[4]
rlabel metal2 103096 2086 103096 2086 0 Q0[5]
rlabel metal2 105784 2086 105784 2086 0 Q0[6]
rlabel metal2 108584 3416 108584 3416 0 Q0[7]
rlabel metal2 111720 2800 111720 2800 0 Q1[0]
rlabel metal2 113848 2086 113848 2086 0 Q1[1]
rlabel metal2 116536 2086 116536 2086 0 Q1[2]
rlabel metal2 119280 3416 119280 3416 0 Q1[3]
rlabel metal2 121912 2086 121912 2086 0 Q1[4]
rlabel metal2 124600 2086 124600 2086 0 Q1[5]
rlabel metal2 126952 2800 126952 2800 0 Q1[6]
rlabel metal2 129976 2086 129976 2086 0 Q1[7]
rlabel metal2 132664 2086 132664 2086 0 Q2[0]
rlabel metal2 135352 2086 135352 2086 0 Q2[1]
rlabel metal2 138376 2800 138376 2800 0 Q2[2]
rlabel metal2 140728 2086 140728 2086 0 Q2[3]
rlabel metal2 143416 2086 143416 2086 0 Q2[4]
rlabel metal2 146272 3416 146272 3416 0 Q2[5]
rlabel metal2 148904 2184 148904 2184 0 Q2[6]
rlabel metal3 154560 3528 154560 3528 0 Q2[7]
rlabel metal2 155064 3472 155064 3472 0 Q3[0]
rlabel metal2 157136 2184 157136 2184 0 Q3[1]
rlabel metal3 159824 3416 159824 3416 0 Q3[2]
rlabel metal2 162232 2058 162232 2058 0 Q3[3]
rlabel metal2 165536 3192 165536 3192 0 Q3[4]
rlabel metal2 167608 2086 167608 2086 0 Q3[5]
rlabel metal2 170296 2086 170296 2086 0 Q3[6]
rlabel metal2 172984 2086 172984 2086 0 Q3[7]
rlabel metal2 175672 2086 175672 2086 0 Q4[0]
rlabel metal2 178360 2086 178360 2086 0 Q4[1]
rlabel metal2 181048 2086 181048 2086 0 Q4[2]
rlabel metal2 184072 2856 184072 2856 0 Q4[3]
rlabel metal2 186424 2086 186424 2086 0 Q4[4]
rlabel metal2 189112 2086 189112 2086 0 Q4[5]
rlabel metal2 191744 3416 191744 3416 0 Q4[6]
rlabel metal2 194488 2086 194488 2086 0 Q4[7]
rlabel metal2 197176 2086 197176 2086 0 Q5[0]
rlabel metal2 199976 3416 199976 3416 0 Q5[1]
rlabel metal2 203112 2800 203112 2800 0 Q5[2]
rlabel metal2 205240 2086 205240 2086 0 Q5[3]
rlabel metal2 207928 2086 207928 2086 0 Q5[4]
rlabel metal2 210672 3416 210672 3416 0 Q5[5]
rlabel metal2 213304 2086 213304 2086 0 Q5[6]
rlabel metal2 215992 2086 215992 2086 0 Q5[7]
rlabel metal2 156184 47642 156184 47642 0 Q6[0]
rlabel metal2 160216 47642 160216 47642 0 Q6[1]
rlabel metal2 164248 47642 164248 47642 0 Q6[2]
rlabel metal2 168728 46480 168728 46480 0 Q6[3]
rlabel metal2 172424 45976 172424 45976 0 Q6[4]
rlabel metal2 176344 47642 176344 47642 0 Q6[5]
rlabel metal2 180320 45976 180320 45976 0 Q6[6]
rlabel metal2 184072 46480 184072 46480 0 Q6[7]
rlabel metal2 188552 45864 188552 45864 0 Q7[0]
rlabel metal2 192472 47642 192472 47642 0 Q7[1]
rlabel metal2 196504 47642 196504 47642 0 Q7[2]
rlabel metal2 200536 47642 200536 47642 0 Q7[3]
rlabel metal2 204568 47642 204568 47642 0 Q7[4]
rlabel metal2 208600 47642 208600 47642 0 Q7[5]
rlabel metal2 212632 47642 212632 47642 0 Q7[6]
rlabel metal2 216664 47642 216664 47642 0 Q7[7]
rlabel metal2 11032 47642 11032 47642 0 WEb_ram
rlabel metal3 138152 45192 138152 45192 0 _000_
rlabel metal2 139664 44968 139664 44968 0 _001_
rlabel metal2 138040 4816 138040 4816 0 _002_
rlabel metal3 150472 10584 150472 10584 0 _003_
rlabel metal2 160104 10024 160104 10024 0 _004_
rlabel metal2 151760 9800 151760 9800 0 _005_
rlabel metal2 153944 7896 153944 7896 0 _006_
rlabel metal2 148848 11368 148848 11368 0 _007_
rlabel metal3 161336 10696 161336 10696 0 _008_
rlabel metal2 138208 6664 138208 6664 0 _009_
rlabel metal2 139496 7168 139496 7168 0 _010_
rlabel metal2 149800 9520 149800 9520 0 _011_
rlabel metal2 152712 3472 152712 3472 0 _012_
rlabel metal2 152488 3696 152488 3696 0 _013_
rlabel metal3 148344 9576 148344 9576 0 _014_
rlabel metal2 156296 5096 156296 5096 0 _015_
rlabel metal2 155008 4872 155008 4872 0 _016_
rlabel metal2 141512 7280 141512 7280 0 _017_
rlabel metal2 150024 8624 150024 8624 0 _018_
rlabel metal2 140168 6216 140168 6216 0 _019_
rlabel metal2 156856 7224 156856 7224 0 _020_
rlabel metal2 157416 5544 157416 5544 0 _021_
rlabel metal2 155736 8120 155736 8120 0 _022_
rlabel metal2 160664 8288 160664 8288 0 _023_
rlabel metal2 161784 6552 161784 6552 0 _024_
rlabel metal3 160776 10584 160776 10584 0 _025_
rlabel metal2 144312 5376 144312 5376 0 _026_
rlabel metal2 140504 4704 140504 4704 0 _027_
rlabel metal2 156296 10976 156296 10976 0 _028_
rlabel metal2 156072 11312 156072 11312 0 _029_
rlabel metal2 144088 7728 144088 7728 0 _030_
rlabel metal2 142968 7616 142968 7616 0 _031_
rlabel metal2 139160 6776 139160 6776 0 _032_
rlabel metal2 139272 5992 139272 5992 0 _033_
rlabel metal2 159320 7168 159320 7168 0 _034_
rlabel metal3 160776 6552 160776 6552 0 _035_
rlabel metal2 154056 5152 154056 5152 0 _036_
rlabel metal2 153944 4760 153944 4760 0 _037_
rlabel metal3 160216 6440 160216 6440 0 _038_
rlabel metal2 153720 5488 153720 5488 0 _039_
rlabel metal2 156856 9016 156856 9016 0 _040_
rlabel metal2 141960 6384 141960 6384 0 _041_
rlabel metal2 134288 5320 134288 5320 0 _042_
rlabel metal2 140952 6552 140952 6552 0 _043_
rlabel metal2 155232 5096 155232 5096 0 _044_
rlabel metal2 155624 5208 155624 5208 0 _045_
rlabel metal2 162904 5264 162904 5264 0 _046_
rlabel metal2 156296 9520 156296 9520 0 _047_
rlabel metal2 156464 5320 156464 5320 0 _048_
rlabel metal3 136136 5320 136136 5320 0 _049_
rlabel metal2 138936 6160 138936 6160 0 _050_
rlabel metal2 151480 6048 151480 6048 0 _051_
rlabel metal2 157416 4424 157416 4424 0 _052_
rlabel metal2 163800 4704 163800 4704 0 _053_
rlabel metal2 157304 5152 157304 5152 0 _054_
rlabel metal2 164360 7336 164360 7336 0 _055_
rlabel metal2 157192 5376 157192 5376 0 _056_
rlabel metal2 156968 11032 156968 11032 0 _057_
rlabel metal2 156744 7112 156744 7112 0 _058_
rlabel metal3 140840 5768 140840 5768 0 _059_
rlabel metal2 130536 6384 130536 6384 0 _060_
rlabel metal2 133224 7840 133224 7840 0 _061_
rlabel metal2 148176 4984 148176 4984 0 _062_
rlabel metal2 146664 4704 146664 4704 0 _063_
rlabel metal2 143304 7840 143304 7840 0 _064_
rlabel metal2 134232 7168 134232 7168 0 _065_
rlabel metal3 150752 5880 150752 5880 0 _066_
rlabel metal2 152264 5488 152264 5488 0 _067_
rlabel metal2 162232 4368 162232 4368 0 _068_
rlabel metal2 162008 4480 162008 4480 0 _069_
rlabel metal2 162456 4200 162456 4200 0 _070_
rlabel metal2 163128 5544 163128 5544 0 _071_
rlabel metal3 164080 4424 164080 4424 0 _072_
rlabel metal2 162568 10136 162568 10136 0 _073_
rlabel metal2 163576 10976 163576 10976 0 _074_
rlabel metal2 163240 4312 163240 4312 0 _075_
rlabel metal2 135128 4368 135128 4368 0 _076_
rlabel metal2 131768 6104 131768 6104 0 _077_
rlabel metal2 135576 8120 135576 8120 0 _078_
rlabel metal2 161896 5488 161896 5488 0 _079_
rlabel metal2 161784 4760 161784 4760 0 _080_
rlabel metal3 163912 5096 163912 5096 0 _081_
rlabel metal2 161112 6048 161112 6048 0 _082_
rlabel metal2 136472 8008 136472 8008 0 _083_
rlabel metal2 131320 5992 131320 5992 0 _084_
rlabel metal3 142520 4816 142520 4816 0 _085_
rlabel metal2 163352 5152 163352 5152 0 _086_
rlabel metal2 163688 6160 163688 6160 0 _087_
rlabel metal2 163800 5320 163800 5320 0 _088_
rlabel metal2 164024 5152 164024 5152 0 _089_
rlabel metal2 139384 4648 139384 4648 0 _090_
rlabel metal2 132104 4984 132104 4984 0 _091_
rlabel metal2 137704 7504 137704 7504 0 _092_
rlabel metal2 163352 6048 163352 6048 0 _093_
rlabel metal2 163240 6608 163240 6608 0 _094_
rlabel metal2 163016 6384 163016 6384 0 _095_
rlabel metal2 162512 5880 162512 5880 0 _096_
rlabel metal2 138488 7784 138488 7784 0 _097_
rlabel metal2 110376 7112 110376 7112 0 _098_
rlabel metal2 137704 9688 137704 9688 0 _099_
rlabel metal2 160776 5712 160776 5712 0 _100_
rlabel metal2 160664 6384 160664 6384 0 _101_
rlabel metal2 160440 6384 160440 6384 0 _102_
rlabel metal2 160216 8120 160216 8120 0 _103_
rlabel metal2 139160 10752 139160 10752 0 _104_
rlabel metal2 136248 43008 136248 43008 0 _105_
rlabel metal2 15064 47642 15064 47642 0 bus_in[0]
rlabel metal2 19096 47642 19096 47642 0 bus_in[1]
rlabel metal2 23128 47642 23128 47642 0 bus_in[2]
rlabel metal2 27832 46200 27832 46200 0 bus_in[3]
rlabel metal2 31640 46480 31640 46480 0 bus_in[4]
rlabel metal2 35504 45976 35504 45976 0 bus_in[5]
rlabel metal2 39256 47642 39256 47642 0 bus_in[6]
rlabel metal2 43232 45976 43232 45976 0 bus_in[7]
rlabel metal2 47768 46760 47768 46760 0 bus_out[0]
rlabel metal2 51800 46312 51800 46312 0 bus_out[1]
rlabel metal2 55384 48174 55384 48174 0 bus_out[2]
rlabel metal2 59752 46760 59752 46760 0 bus_out[3]
rlabel metal2 63504 46088 63504 46088 0 bus_out[4]
rlabel metal2 67480 47642 67480 47642 0 bus_out[5]
rlabel metal2 71512 47642 71512 47642 0 bus_out[6]
rlabel metal2 75544 47138 75544 47138 0 bus_out[7]
rlabel metal2 124264 36680 124264 36680 0 clknet_0_wb_clk_i
rlabel metal2 101304 29904 101304 29904 0 clknet_1_0__leaf_wb_clk_i
rlabel metal2 125384 29904 125384 29904 0 clknet_1_1__leaf_wb_clk_i
rlabel metal2 116872 4480 116872 4480 0 net1
rlabel metal2 114464 3416 114464 3416 0 net10
rlabel metal2 52024 4368 52024 4368 0 net100
rlabel metal2 5656 4592 5656 4592 0 net101
rlabel metal2 50456 4200 50456 4200 0 net102
rlabel metal2 53144 4200 53144 4200 0 net103
rlabel metal2 55832 4592 55832 4592 0 net104
rlabel metal2 58520 4200 58520 4200 0 net105
rlabel metal2 61208 4200 61208 4200 0 net106
rlabel metal2 63896 4200 63896 4200 0 net107
rlabel metal2 66584 4592 66584 4592 0 net108
rlabel metal2 69272 4200 69272 4200 0 net109
rlabel metal2 117096 3584 117096 3584 0 net11
rlabel metal2 77224 4032 77224 4032 0 net110
rlabel metal2 80584 3304 80584 3304 0 net111
rlabel metal3 82824 4312 82824 4312 0 net112
rlabel metal3 86184 3416 86184 3416 0 net113
rlabel metal3 87584 4312 87584 4312 0 net114
rlabel metal2 89040 4536 89040 4536 0 net115
rlabel metal2 152824 45752 152824 45752 0 net116
rlabel metal2 140952 9184 140952 9184 0 net117
rlabel metal3 51744 45640 51744 45640 0 net118
rlabel metal3 54656 45864 54656 45864 0 net119
rlabel metal2 120120 3808 120120 3808 0 net12
rlabel metal2 138040 10192 138040 10192 0 net120
rlabel metal2 69720 30800 69720 30800 0 net121
rlabel metal2 65912 45808 65912 45808 0 net122
rlabel metal3 71848 45640 71848 45640 0 net123
rlabel metal3 75320 45640 75320 45640 0 net124
rlabel metal2 78624 45080 78624 45080 0 net125
rlabel metal2 6328 2030 6328 2030 0 net126
rlabel metal2 9016 2030 9016 2030 0 net127
rlabel metal2 11704 2030 11704 2030 0 net128
rlabel metal2 14392 2030 14392 2030 0 net129
rlabel metal2 122472 2856 122472 2856 0 net13
rlabel metal2 17080 2030 17080 2030 0 net130
rlabel metal2 19768 854 19768 854 0 net131
rlabel metal2 22456 2030 22456 2030 0 net132
rlabel metal2 25144 2030 25144 2030 0 net133
rlabel metal2 125160 4704 125160 4704 0 net14
rlabel metal4 137816 4536 137816 4536 0 net15
rlabel metal3 143416 4592 143416 4592 0 net16
rlabel metal2 133224 3864 133224 3864 0 net17
rlabel metal2 138936 5040 138936 5040 0 net18
rlabel metal2 139160 4200 139160 4200 0 net19
rlabel metal2 93464 3864 93464 3864 0 net2
rlabel metal2 141288 3864 141288 3864 0 net20
rlabel metal2 143976 4648 143976 4648 0 net21
rlabel metal2 146776 4256 146776 4256 0 net22
rlabel metal2 149352 5432 149352 5432 0 net23
rlabel metal2 153048 4032 153048 4032 0 net24
rlabel metal2 155288 3640 155288 3640 0 net25
rlabel metal2 157864 4144 157864 4144 0 net26
rlabel metal3 158928 4872 158928 4872 0 net27
rlabel metal2 163352 3640 163352 3640 0 net28
rlabel metal2 165480 3864 165480 3864 0 net29
rlabel metal2 95592 3528 95592 3528 0 net3
rlabel metal3 165592 6776 165592 6776 0 net30
rlabel metal2 170520 5320 170520 5320 0 net31
rlabel metal2 173208 3584 173208 3584 0 net32
rlabel metal2 175896 3584 175896 3584 0 net33
rlabel metal2 178584 4144 178584 4144 0 net34
rlabel metal2 181272 4592 181272 4592 0 net35
rlabel metal2 184520 3752 184520 3752 0 net36
rlabel metal2 186648 3528 186648 3528 0 net37
rlabel metal2 189336 4704 189336 4704 0 net38
rlabel metal2 192136 4648 192136 4648 0 net39
rlabel metal2 98280 4032 98280 4032 0 net4
rlabel metal2 194712 4480 194712 4480 0 net40
rlabel metal2 140280 4256 140280 4256 0 net41
rlabel metal2 141848 5264 141848 5264 0 net42
rlabel metal2 144368 6440 144368 6440 0 net43
rlabel metal2 206024 3416 206024 3416 0 net44
rlabel metal2 208712 2464 208712 2464 0 net45
rlabel metal3 196560 3584 196560 3584 0 net46
rlabel metal2 213976 5264 213976 5264 0 net47
rlabel metal2 216664 4088 216664 4088 0 net48
rlabel metal2 156744 44660 156744 44660 0 net49
rlabel metal2 101080 3472 101080 3472 0 net5
rlabel metal2 157192 9632 157192 9632 0 net50
rlabel metal2 157752 11536 157752 11536 0 net51
rlabel metal2 169288 29904 169288 29904 0 net52
rlabel metal2 173096 44688 173096 44688 0 net53
rlabel metal2 176904 28840 176904 28840 0 net54
rlabel metal2 168056 13048 168056 13048 0 net55
rlabel metal3 173768 15960 173768 15960 0 net56
rlabel metal3 143248 3640 143248 3640 0 net57
rlabel metal2 142520 5152 142520 5152 0 net58
rlabel metal3 171584 17640 171584 17640 0 net59
rlabel metal2 103656 3752 103656 3752 0 net6
rlabel metal3 165312 2408 165312 2408 0 net60
rlabel metal3 177800 45976 177800 45976 0 net61
rlabel metal2 209384 30016 209384 30016 0 net62
rlabel metal2 213976 29232 213976 29232 0 net63
rlabel metal3 211680 45976 211680 45976 0 net64
rlabel metal3 138992 44968 138992 44968 0 net65
rlabel metal2 49784 6384 49784 6384 0 net66
rlabel metal2 52472 5096 52472 5096 0 net67
rlabel metal2 23912 35952 23912 35952 0 net68
rlabel metal2 28952 29288 28952 29288 0 net69
rlabel metal2 106512 3416 106512 3416 0 net7
rlabel metal3 37800 45416 37800 45416 0 net70
rlabel metal3 37184 45864 37184 45864 0 net71
rlabel metal2 65856 5208 65856 5208 0 net72
rlabel metal3 46032 45864 46032 45864 0 net73
rlabel metal2 80136 44632 80136 44632 0 net74
rlabel metal3 133168 30072 133168 30072 0 net75
rlabel metal2 122024 5208 122024 5208 0 net76
rlabel metal2 126392 5208 126392 5208 0 net77
rlabel metal2 132664 45024 132664 45024 0 net78
rlabel metal2 135912 44912 135912 44912 0 net79
rlabel metal2 109032 4256 109032 4256 0 net8
rlabel metal2 140280 44660 140280 44660 0 net80
rlabel metal2 139832 44408 139832 44408 0 net81
rlabel metal2 135800 29568 135800 29568 0 net82
rlabel metal2 92232 43400 92232 43400 0 net83
rlabel metal2 93352 5152 93352 5152 0 net84
rlabel metal2 98168 5208 98168 5208 0 net85
rlabel metal2 101864 5208 101864 5208 0 net86
rlabel metal2 106120 5152 106120 5152 0 net87
rlabel metal2 109704 5152 109704 5152 0 net88
rlabel metal2 116704 31192 116704 31192 0 net89
rlabel metal2 112560 3416 112560 3416 0 net9
rlabel metal2 118104 5152 118104 5152 0 net90
rlabel metal3 6832 5208 6832 5208 0 net91
rlabel metal2 31528 4704 31528 4704 0 net92
rlabel metal2 97496 6048 97496 6048 0 net93
rlabel metal2 101080 4760 101080 4760 0 net94
rlabel metal2 39256 5208 39256 5208 0 net95
rlabel metal2 94024 4424 94024 4424 0 net96
rlabel metal2 44520 5264 44520 5264 0 net97
rlabel metal2 46984 4704 46984 4704 0 net98
rlabel metal2 50568 3920 50568 3920 0 net99
rlabel metal2 79576 47642 79576 47642 0 ram_enabled
rlabel metal2 83608 47642 83608 47642 0 requested_addr[0]
rlabel metal2 123928 47642 123928 47642 0 requested_addr[10]
rlabel metal2 127960 47642 127960 47642 0 requested_addr[11]
rlabel metal2 131992 47642 131992 47642 0 requested_addr[12]
rlabel metal2 136024 47642 136024 47642 0 requested_addr[13]
rlabel metal2 140056 47642 140056 47642 0 requested_addr[14]
rlabel metal2 144088 47642 144088 47642 0 requested_addr[15]
rlabel metal2 87640 47642 87640 47642 0 requested_addr[1]
rlabel metal2 91672 47642 91672 47642 0 requested_addr[2]
rlabel metal2 95704 47642 95704 47642 0 requested_addr[3]
rlabel metal2 100184 46480 100184 46480 0 requested_addr[4]
rlabel metal2 103880 45976 103880 45976 0 requested_addr[5]
rlabel metal2 107800 47642 107800 47642 0 requested_addr[6]
rlabel metal2 111776 45976 111776 45976 0 requested_addr[7]
rlabel metal2 115528 46424 115528 46424 0 requested_addr[8]
rlabel metal2 120008 45864 120008 45864 0 requested_addr[9]
rlabel metal2 135856 30296 135856 30296 0 requested_addr_latch\[0\]
rlabel metal2 134792 43568 134792 43568 0 requested_addr_latch\[12\]
rlabel metal2 138040 44044 138040 44044 0 requested_addr_latch\[13\]
rlabel metal2 137592 43176 137592 43176 0 requested_addr_latch\[14\]
rlabel metal2 141624 44744 141624 44744 0 requested_addr_latch\[15\]
rlabel metal2 137928 20384 137928 20384 0 requested_addr_latch\[1\]
rlabel metal2 140280 22176 140280 22176 0 requested_addr_latch\[2\]
rlabel metal2 7000 47642 7000 47642 0 rst
rlabel metal2 2968 43218 2968 43218 0 wb_clk_i
<< properties >>
string FIXED_BBOX 0 0 220000 50000
<< end >>
