VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO boot_rom
  CLASS BLOCK ;
  FOREIGN boot_rom ;
  ORIGIN 0.000 0.000 ;
  SIZE 210.000 BY 210.000 ;
  PIN bus_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 79.520 206.000 80.080 210.000 ;
    END
  END bus_out[0]
  PIN bus_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 96.320 206.000 96.880 210.000 ;
    END
  END bus_out[1]
  PIN bus_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 113.120 206.000 113.680 210.000 ;
    END
  END bus_out[2]
  PIN bus_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 129.920 206.000 130.480 210.000 ;
    END
  END bus_out[3]
  PIN bus_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 146.720 206.000 147.280 210.000 ;
    END
  END bus_out[4]
  PIN bus_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 163.520 206.000 164.080 210.000 ;
    END
  END bus_out[5]
  PIN bus_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 180.320 206.000 180.880 210.000 ;
    END
  END bus_out[6]
  PIN bus_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 197.120 206.000 197.680 210.000 ;
    END
  END bus_out[7]
  PIN cs_port[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 29.120 206.000 29.680 210.000 ;
    END
  END cs_port[0]
  PIN cs_port[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 45.920 206.000 46.480 210.000 ;
    END
  END cs_port[1]
  PIN cs_port[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 62.720 206.000 63.280 210.000 ;
    END
  END cs_port[2]
  PIN last_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 160.160 4.000 160.720 ;
    END
  END last_addr[0]
  PIN last_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 164.640 4.000 165.200 ;
    END
  END last_addr[1]
  PIN last_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 169.120 4.000 169.680 ;
    END
  END last_addr[2]
  PIN last_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 173.600 4.000 174.160 ;
    END
  END last_addr[3]
  PIN last_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 178.080 4.000 178.640 ;
    END
  END last_addr[4]
  PIN last_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 182.560 4.000 183.120 ;
    END
  END last_addr[5]
  PIN last_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 187.040 4.000 187.600 ;
    END
  END last_addr[6]
  PIN last_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 191.520 4.000 192.080 ;
    END
  END last_addr[7]
  PIN ram_end[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 88.480 4.000 89.040 ;
    END
  END ram_end[0]
  PIN ram_end[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 133.280 4.000 133.840 ;
    END
  END ram_end[10]
  PIN ram_end[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 137.760 4.000 138.320 ;
    END
  END ram_end[11]
  PIN ram_end[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 142.240 4.000 142.800 ;
    END
  END ram_end[12]
  PIN ram_end[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 146.720 4.000 147.280 ;
    END
  END ram_end[13]
  PIN ram_end[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 151.200 4.000 151.760 ;
    END
  END ram_end[14]
  PIN ram_end[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 155.680 4.000 156.240 ;
    END
  END ram_end[15]
  PIN ram_end[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 92.960 4.000 93.520 ;
    END
  END ram_end[1]
  PIN ram_end[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 97.440 4.000 98.000 ;
    END
  END ram_end[2]
  PIN ram_end[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 101.920 4.000 102.480 ;
    END
  END ram_end[3]
  PIN ram_end[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 106.400 4.000 106.960 ;
    END
  END ram_end[4]
  PIN ram_end[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 110.880 4.000 111.440 ;
    END
  END ram_end[5]
  PIN ram_end[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 115.360 4.000 115.920 ;
    END
  END ram_end[6]
  PIN ram_end[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 119.840 4.000 120.400 ;
    END
  END ram_end[7]
  PIN ram_end[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 124.320 4.000 124.880 ;
    END
  END ram_end[8]
  PIN ram_end[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 128.800 4.000 129.360 ;
    END
  END ram_end[9]
  PIN ram_start[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 16.800 4.000 17.360 ;
    END
  END ram_start[0]
  PIN ram_start[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 61.600 4.000 62.160 ;
    END
  END ram_start[10]
  PIN ram_start[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 66.080 4.000 66.640 ;
    END
  END ram_start[11]
  PIN ram_start[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 70.560 4.000 71.120 ;
    END
  END ram_start[12]
  PIN ram_start[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 75.040 4.000 75.600 ;
    END
  END ram_start[13]
  PIN ram_start[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 79.520 4.000 80.080 ;
    END
  END ram_start[14]
  PIN ram_start[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 84.000 4.000 84.560 ;
    END
  END ram_start[15]
  PIN ram_start[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 21.280 4.000 21.840 ;
    END
  END ram_start[1]
  PIN ram_start[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 25.760 4.000 26.320 ;
    END
  END ram_start[2]
  PIN ram_start[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 30.240 4.000 30.800 ;
    END
  END ram_start[3]
  PIN ram_start[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 34.720 4.000 35.280 ;
    END
  END ram_start[4]
  PIN ram_start[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 39.200 4.000 39.760 ;
    END
  END ram_start[5]
  PIN ram_start[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 43.680 4.000 44.240 ;
    END
  END ram_start[6]
  PIN ram_start[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 48.160 4.000 48.720 ;
    END
  END ram_start[7]
  PIN ram_start[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 52.640 4.000 53.200 ;
    END
  END ram_start[8]
  PIN ram_start[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 57.120 4.000 57.680 ;
    END
  END ram_start[9]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 192.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 192.380 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 192.380 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 12.320 206.000 12.880 210.000 ;
    END
  END wb_clk_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 203.280 193.050 ;
      LAYER Metal2 ;
        RECT 5.740 205.700 12.020 206.500 ;
        RECT 13.180 205.700 28.820 206.500 ;
        RECT 29.980 205.700 45.620 206.500 ;
        RECT 46.780 205.700 62.420 206.500 ;
        RECT 63.580 205.700 79.220 206.500 ;
        RECT 80.380 205.700 96.020 206.500 ;
        RECT 97.180 205.700 112.820 206.500 ;
        RECT 113.980 205.700 129.620 206.500 ;
        RECT 130.780 205.700 146.420 206.500 ;
        RECT 147.580 205.700 163.220 206.500 ;
        RECT 164.380 205.700 180.020 206.500 ;
        RECT 181.180 205.700 196.820 206.500 ;
        RECT 5.740 15.490 197.540 205.700 ;
      LAYER Metal3 ;
        RECT 4.300 191.220 188.630 192.220 ;
        RECT 4.000 187.900 188.630 191.220 ;
        RECT 4.300 186.740 188.630 187.900 ;
        RECT 4.000 183.420 188.630 186.740 ;
        RECT 4.300 182.260 188.630 183.420 ;
        RECT 4.000 178.940 188.630 182.260 ;
        RECT 4.300 177.780 188.630 178.940 ;
        RECT 4.000 174.460 188.630 177.780 ;
        RECT 4.300 173.300 188.630 174.460 ;
        RECT 4.000 169.980 188.630 173.300 ;
        RECT 4.300 168.820 188.630 169.980 ;
        RECT 4.000 165.500 188.630 168.820 ;
        RECT 4.300 164.340 188.630 165.500 ;
        RECT 4.000 161.020 188.630 164.340 ;
        RECT 4.300 159.860 188.630 161.020 ;
        RECT 4.000 156.540 188.630 159.860 ;
        RECT 4.300 155.380 188.630 156.540 ;
        RECT 4.000 152.060 188.630 155.380 ;
        RECT 4.300 150.900 188.630 152.060 ;
        RECT 4.000 147.580 188.630 150.900 ;
        RECT 4.300 146.420 188.630 147.580 ;
        RECT 4.000 143.100 188.630 146.420 ;
        RECT 4.300 141.940 188.630 143.100 ;
        RECT 4.000 138.620 188.630 141.940 ;
        RECT 4.300 137.460 188.630 138.620 ;
        RECT 4.000 134.140 188.630 137.460 ;
        RECT 4.300 132.980 188.630 134.140 ;
        RECT 4.000 129.660 188.630 132.980 ;
        RECT 4.300 128.500 188.630 129.660 ;
        RECT 4.000 125.180 188.630 128.500 ;
        RECT 4.300 124.020 188.630 125.180 ;
        RECT 4.000 120.700 188.630 124.020 ;
        RECT 4.300 119.540 188.630 120.700 ;
        RECT 4.000 116.220 188.630 119.540 ;
        RECT 4.300 115.060 188.630 116.220 ;
        RECT 4.000 111.740 188.630 115.060 ;
        RECT 4.300 110.580 188.630 111.740 ;
        RECT 4.000 107.260 188.630 110.580 ;
        RECT 4.300 106.100 188.630 107.260 ;
        RECT 4.000 102.780 188.630 106.100 ;
        RECT 4.300 101.620 188.630 102.780 ;
        RECT 4.000 98.300 188.630 101.620 ;
        RECT 4.300 97.140 188.630 98.300 ;
        RECT 4.000 93.820 188.630 97.140 ;
        RECT 4.300 92.660 188.630 93.820 ;
        RECT 4.000 89.340 188.630 92.660 ;
        RECT 4.300 88.180 188.630 89.340 ;
        RECT 4.000 84.860 188.630 88.180 ;
        RECT 4.300 83.700 188.630 84.860 ;
        RECT 4.000 80.380 188.630 83.700 ;
        RECT 4.300 79.220 188.630 80.380 ;
        RECT 4.000 75.900 188.630 79.220 ;
        RECT 4.300 74.740 188.630 75.900 ;
        RECT 4.000 71.420 188.630 74.740 ;
        RECT 4.300 70.260 188.630 71.420 ;
        RECT 4.000 66.940 188.630 70.260 ;
        RECT 4.300 65.780 188.630 66.940 ;
        RECT 4.000 62.460 188.630 65.780 ;
        RECT 4.300 61.300 188.630 62.460 ;
        RECT 4.000 57.980 188.630 61.300 ;
        RECT 4.300 56.820 188.630 57.980 ;
        RECT 4.000 53.500 188.630 56.820 ;
        RECT 4.300 52.340 188.630 53.500 ;
        RECT 4.000 49.020 188.630 52.340 ;
        RECT 4.300 47.860 188.630 49.020 ;
        RECT 4.000 44.540 188.630 47.860 ;
        RECT 4.300 43.380 188.630 44.540 ;
        RECT 4.000 40.060 188.630 43.380 ;
        RECT 4.300 38.900 188.630 40.060 ;
        RECT 4.000 35.580 188.630 38.900 ;
        RECT 4.300 34.420 188.630 35.580 ;
        RECT 4.000 31.100 188.630 34.420 ;
        RECT 4.300 29.940 188.630 31.100 ;
        RECT 4.000 26.620 188.630 29.940 ;
        RECT 4.300 25.460 188.630 26.620 ;
        RECT 4.000 22.140 188.630 25.460 ;
        RECT 4.300 20.980 188.630 22.140 ;
        RECT 4.000 17.660 188.630 20.980 ;
        RECT 4.300 16.500 188.630 17.660 ;
        RECT 4.000 15.540 188.630 16.500 ;
      LAYER Metal4 ;
        RECT 11.900 40.410 21.940 189.750 ;
        RECT 24.140 40.410 98.740 189.750 ;
        RECT 100.940 40.410 121.380 189.750 ;
  END
END boot_rom
END LIBRARY

