// This is the unpowered netlist.
module boot_rom (WEb_raw,
    le_hi_act,
    le_lo_act,
    rom_enabled,
    rst,
    wb_clk_i,
    bus_in,
    bus_out,
    cs_port,
    ram_end,
    ram_start);
 input WEb_raw;
 input le_hi_act;
 input le_lo_act;
 input rom_enabled;
 input rst;
 input wb_clk_i;
 input [7:0] bus_in;
 output [7:0] bus_out;
 input [2:0] cs_port;
 input [15:0] ram_end;
 input [15:0] ram_start;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire clknet_0_wb_clk_i;
 wire clknet_2_0__leaf_wb_clk_i;
 wire clknet_2_1__leaf_wb_clk_i;
 wire clknet_2_2__leaf_wb_clk_i;
 wire clknet_2_3__leaf_wb_clk_i;
 wire \full_addr[0] ;
 wire \full_addr[10] ;
 wire \full_addr[11] ;
 wire \full_addr[12] ;
 wire \full_addr[13] ;
 wire \full_addr[14] ;
 wire \full_addr[15] ;
 wire \full_addr[1] ;
 wire \full_addr[2] ;
 wire \full_addr[3] ;
 wire \full_addr[4] ;
 wire \full_addr[5] ;
 wire \full_addr[6] ;
 wire \full_addr[7] ;
 wire \full_addr[8] ;
 wire \full_addr[9] ;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire \writable[0] ;
 wire \writable[10] ;
 wire \writable[11] ;
 wire \writable[12] ;
 wire \writable[13] ;
 wire \writable[14] ;
 wire \writable[15] ;
 wire \writable[1] ;
 wire \writable[2] ;
 wire \writable[3] ;
 wire \writable[4] ;
 wire \writable[5] ;
 wire \writable[6] ;
 wire \writable[7] ;
 wire \writable[8] ;
 wire \writable[9] ;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0567__I (.I(\full_addr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0584__A1 (.I(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0584__A2 (.I(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0585__I (.I(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0586__I (.I(\full_addr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0612__A3 (.I(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0619__I (.I(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0622__I (.I(\full_addr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0636__A3 (.I(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0636__B1 (.I(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0637__A1 (.I(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0637__B1 (.I(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0637__B2 (.I(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0644__A1 (.I(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0644__A2 (.I(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0647__I (.I(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0653__A1 (.I(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0653__B1 (.I(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0653__B2 (.I(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0657__I (.I(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0659__A1 (.I(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0659__A2 (.I(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0659__B (.I(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0665__A2 (.I(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0668__I (.I(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0669__A1 (.I(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0674__I (.I(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0675__A1 (.I(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0675__A2 (.I(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0677__I (.I(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0679__A1 (.I(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0680__I (.I(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0681__A1 (.I(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0683__A2 (.I(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0686__I (.I(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0692__B2 (.I(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0693__A1 (.I(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0693__A2 (.I(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0699__B (.I(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0700__A3 (.I(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0701__A1 (.I(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0701__A2 (.I(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0704__I (.I(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0706__A2 (.I(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0708__A1 (.I(\full_addr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0709__I (.I(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0716__I (.I(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0718__A2 (.I(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0718__B1 (.I(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0719__A1 (.I(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0723__I (.I(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0726__A3 (.I(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0727__I (.I(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0729__A2 (.I(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0733__A2 (.I(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0733__B1 (.I(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0733__B2 (.I(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0735__A1 (.I(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0737__A4 (.I(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0743__A3 (.I(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0743__B2 (.I(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0744__A1 (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0744__C (.I(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0745__A2 (.I(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0747__A1 (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0747__A2 (.I(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0748__A3 (.I(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0752__I (.I(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0755__I (.I(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0756__A2 (.I(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0756__B (.I(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0759__I (.I(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0761__A3 (.I(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0763__I (.I(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0765__A1 (.I(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0765__A2 (.I(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0768__I (.I(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0769__A1 (.I(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0769__A2 (.I(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0771__A1 (.I(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0771__A2 (.I(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0771__B (.I(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0774__I (.I(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0777__A1 (.I(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0777__A2 (.I(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0777__B2 (.I(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0778__I (.I(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0779__A1 (.I(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0779__B2 (.I(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0779__C1 (.I(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0779__C2 (.I(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0780__A3 (.I(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0783__A1 (.I(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0783__A2 (.I(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0783__B1 (.I(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0783__B2 (.I(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0783__C2 (.I(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0786__A1 (.I(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0786__A2 (.I(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0786__B (.I(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0788__B1 (.I(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0788__B2 (.I(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0788__C1 (.I(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0788__C2 (.I(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0793__A1 (.I(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0793__A2 (.I(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0793__B1 (.I(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0793__C1 (.I(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0793__C2 (.I(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0795__A1 (.I(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0798__I (.I(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0799__A2 (.I(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0800__I (.I(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0801__A1 (.I(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0802__B (.I(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0805__A2 (.I(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0809__A1 (.I(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0809__B (.I(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0811__I (.I(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0812__A2 (.I(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0812__A3 (.I(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0815__A2 (.I(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0816__A1 (.I(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0818__A1 (.I(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0818__A2 (.I(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0819__A1 (.I(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0819__A2 (.I(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0820__A1 (.I(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0820__A2 (.I(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0821__B (.I(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0821__C (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0826__A2 (.I(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0827__A2 (.I(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0827__B1 (.I(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0832__A1 (.I(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0833__C1 (.I(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0833__C2 (.I(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0834__I (.I(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0835__A1 (.I(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0836__A1 (.I(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0837__I (.I(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0842__A2 (.I(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0843__A1 (.I(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0843__A2 (.I(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0847__A2 (.I(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0848__B1 (.I(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0848__B2 (.I(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0850__A1 (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0850__A2 (.I(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0851__A2 (.I(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0852__A2 (.I(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0852__B2 (.I(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0859__A1 (.I(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0859__A2 (.I(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0860__A1 (.I(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0860__A2 (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0861__A1 (.I(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0861__A2 (.I(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0861__B (.I(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0862__A1 (.I(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0862__B1 (.I(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0862__B2 (.I(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0864__A1 (.I(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0866__B2 (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0868__A1 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0870__A1 (.I(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0870__A2 (.I(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0870__B1 (.I(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0872__I (.I(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0875__A1 (.I(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0876__I (.I(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0877__A1 (.I(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0877__A2 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0878__I (.I(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0880__A1 (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0881__I (.I(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0883__B1 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0883__B2 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0893__A2 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0894__A1 (.I(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0894__A2 (.I(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0896__A1 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0897__A2 (.I(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0898__B1 (.I(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0899__A2 (.I(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0899__B (.I(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0903__A1 (.I(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0903__A2 (.I(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0905__A1 (.I(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0905__C1 (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0906__A2 (.I(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0907__A1 (.I(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0907__A2 (.I(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0908__A1 (.I(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0908__B1 (.I(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0910__A2 (.I(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0910__A3 (.I(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0910__A4 (.I(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0914__A1 (.I(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0919__A1 (.I(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0919__A2 (.I(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0920__A1 (.I(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0921__A2 (.I(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0922__A1 (.I(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0923__A1 (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0924__A1 (.I(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0924__A2 (.I(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0928__A1 (.I(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0928__A2 (.I(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0929__A1 (.I(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0930__B1 (.I(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0930__B2 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0931__A1 (.I(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0932__A2 (.I(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0934__A2 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0937__I (.I(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0938__I (.I(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0939__A2 (.I(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0939__B (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0940__A1 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0940__B (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0941__A1 (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0942__A1 (.I(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0950__A3 (.I(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0953__I (.I(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0954__A2 (.I(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0955__A1 (.I(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0955__A2 (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0957__A1 (.I(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0957__B (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0959__B2 (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0960__A1 (.I(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0961__A1 (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0961__A3 (.I(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0967__A1 (.I(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0974__A1 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0974__A2 (.I(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0976__A2 (.I(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0977__A1 (.I(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0979__A2 (.I(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0980__A1 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0980__A2 (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0980__B1 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0981__A1 (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0981__C2 (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0983__A4 (.I(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0986__A1 (.I(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0987__A1 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0988__A3 (.I(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0989__A1 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0989__B (.I(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0990__A1 (.I(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0991__B1 (.I(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0991__B2 (.I(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0992__A1 (.I(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0994__A1 (.I(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0995__A3 (.I(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0998__B (.I(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__0998__C (.I(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1001__A1 (.I(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1002__A3 (.I(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1003__A1 (.I(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1003__A2 (.I(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1003__B2 (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1005__A1 (.I(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1009__A1 (.I(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1012__A1 (.I(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1012__A3 (.I(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1012__A4 (.I(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1013__C2 (.I(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1014__A3 (.I(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1017__A1 (.I(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1021__A1 (.I(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1023__A1 (.I(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1024__A1 (.I(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1031__A1 (.I(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1034__I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1037__I (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1038__I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1039__A1 (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1040__A1 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1042__A1 (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1043__A1 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1045__A1 (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1046__A1 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1048__I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1049__A1 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1050__A1 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1052__I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1053__I (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1054__A1 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1055__A1 (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1057__A1 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1058__A1 (.I(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1060__A1 (.I(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1061__A1 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1063__A2 (.I(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1064__A1 (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1065__A2 (.I(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1066__I (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1067__I (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1069__I (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1071__A1 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1073__A1 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1075__A1 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1077__A1 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1078__I (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1079__I (.I(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1080__I (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1082__A1 (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1084__A1 (.I(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1086__A1 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1088__A1 (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1089__I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1090__I (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1091__I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1093__A1 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1095__A1 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1097__A1 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1098__I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1100__A1 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1101__I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1102__I (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1104__A1 (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1106__A1 (.I(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1108__A1 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1110__A1 (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1114__I (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1116__A1 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1118__A1 (.I(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1120__A1 (.I(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1122__A1 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1125__I (.I(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1127__A1 (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1129__A1 (.I(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1131__A1 (.I(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1133__A1 (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1134__CLK (.I(clknet_2_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1135__CLK (.I(clknet_2_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1136__CLK (.I(clknet_2_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1137__CLK (.I(clknet_2_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1146__CLK (.I(clknet_2_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1150__CLK (.I(clknet_2_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1152__CLK (.I(clknet_2_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1153__CLK (.I(clknet_2_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1154__CLK (.I(clknet_2_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1155__CLK (.I(clknet_2_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1156__CLK (.I(clknet_2_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1157__CLK (.I(clknet_2_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1158__CLK (.I(clknet_2_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1159__CLK (.I(clknet_2_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1160__CLK (.I(clknet_2_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1162__CLK (.I(clknet_2_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1163__CLK (.I(clknet_2_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__1165__CLK (.I(clknet_2_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_wb_clk_i_I (.I(wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_0__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_1__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_2__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_2_3__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(cs_port[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(cs_port[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(cs_port[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(le_hi_act));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(le_lo_act));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(ram_end[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(ram_end[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(ram_end[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(ram_end[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(ram_end[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(WEb_raw));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(ram_end[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(ram_end[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(ram_end[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(ram_end[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(ram_end[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(ram_end[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(ram_end[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(ram_end[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(ram_end[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(ram_end[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(bus_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(ram_end[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(ram_start[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(ram_start[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(ram_start[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input34_I (.I(ram_start[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input35_I (.I(ram_start[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input36_I (.I(ram_start[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input37_I (.I(ram_start[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input38_I (.I(ram_start[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input39_I (.I(ram_start[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(bus_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input40_I (.I(ram_start[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input41_I (.I(ram_start[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input42_I (.I(ram_start[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input43_I (.I(ram_start[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input44_I (.I(ram_start[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input45_I (.I(ram_start[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input46_I (.I(ram_start[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input47_I (.I(rom_enabled));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input48_I (.I(rst));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(bus_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(bus_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(bus_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(bus_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(bus_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(bus_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output49_I (.I(net49));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output50_I (.I(net50));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output51_I (.I(net51));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output52_I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output53_I (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output54_I (.I(net54));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output55_I (.I(net55));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output56_I (.I(net56));
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_0_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_0_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_15_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_16_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_19_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_1_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_20_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_21_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_22_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_25_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_26_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_27_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_28_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_30_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_32_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_34_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_35_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_38_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_40_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_42_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_44_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_46_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_50_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_51_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_52_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_52_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_52_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_53_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_54_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_54_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_54_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_55_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_55_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_55_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_55_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_55_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_55_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_55_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_56_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_56_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_56_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_56_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_56_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_56_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_56_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_57_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_57_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_57_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_57_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_57_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_57_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_58_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_58_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_58_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_58_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_58_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_58_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_59_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_59_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_59_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_59_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_59_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_59_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_59_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_60_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_60_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_60_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_60_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_60_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_60_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_61_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_61_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_61_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_61_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_61_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_61_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_61_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_62_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_62_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_62_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_62_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_62_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_62_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_62_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_63_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_63_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_63_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_63_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_63_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_63_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_64_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_64_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_64_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_64_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_64_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_64_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_64_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_65_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_65_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_65_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_65_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_65_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_65_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_66_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_66_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_66_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_66_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_66_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_67_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_67_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_67_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_67_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Left_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Left_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Left_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Left_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Left_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Left_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Left_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Left_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Left_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Left_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Left_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_55_Right_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Left_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_56_Right_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Left_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_57_Right_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Left_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_58_Right_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Left_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_59_Right_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Left_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_60_Right_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Left_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_61_Right_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Left_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_62_Right_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Left_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_63_Right_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Left_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_64_Right_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Left_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_65_Right_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Left_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_66_Right_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Left_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_67_Right_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_55_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_56_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_57_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_58_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_59_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_60_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_61_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_62_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_63_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_64_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_65_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_66_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_67_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0563_ (.I(\writable[0] ),
    .ZN(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _0564_ (.A1(\full_addr[11] ),
    .A2(\full_addr[10] ),
    .A3(\full_addr[9] ),
    .A4(\full_addr[8] ),
    .Z(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _0565_ (.A1(\full_addr[15] ),
    .A2(\full_addr[14] ),
    .A3(\full_addr[13] ),
    .ZN(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _0566_ (.A1(\full_addr[12] ),
    .A2(_0033_),
    .A3(_0034_),
    .ZN(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _0567_ (.I(\full_addr[7] ),
    .Z(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0568_ (.I(\full_addr[6] ),
    .Z(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _0569_ (.I(_0037_),
    .Z(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0570_ (.I(\full_addr[5] ),
    .Z(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _0571_ (.I(_0039_),
    .Z(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _0572_ (.I(\full_addr[4] ),
    .Z(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _0573_ (.A1(_0036_),
    .A2(_0038_),
    .A3(_0040_),
    .A4(_0041_),
    .ZN(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0574_ (.I(\full_addr[3] ),
    .Z(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0575_ (.I(_0043_),
    .Z(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0576_ (.I(\full_addr[2] ),
    .Z(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0577_ (.I(_0045_),
    .Z(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0578_ (.I(\full_addr[1] ),
    .Z(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0579_ (.I(_0047_),
    .Z(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0580_ (.I(\full_addr[0] ),
    .Z(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0581_ (.I(_0049_),
    .ZN(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0582_ (.I(_0050_),
    .Z(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _0583_ (.A1(_0044_),
    .A2(_0046_),
    .A3(_0048_),
    .A4(_0051_),
    .ZN(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _0584_ (.A1(_0035_),
    .A2(_0042_),
    .A3(_0052_),
    .ZN(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _0585_ (.I(_0053_),
    .Z(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0586_ (.I(\full_addr[7] ),
    .Z(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0587_ (.I(_0055_),
    .Z(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _0588_ (.I(\full_addr[6] ),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _0589_ (.I(_0057_),
    .Z(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _0590_ (.I(_0039_),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0591_ (.I(\full_addr[4] ),
    .Z(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0592_ (.I(_0060_),
    .Z(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _0593_ (.A1(_0056_),
    .A2(_0058_),
    .A3(_0059_),
    .A4(_0061_),
    .ZN(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _0594_ (.I(_0062_),
    .Z(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0595_ (.I(\full_addr[1] ),
    .ZN(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0596_ (.I(_0064_),
    .Z(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0597_ (.I(_0049_),
    .Z(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0598_ (.A1(_0043_),
    .A2(_0045_),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0599_ (.I(_0067_),
    .Z(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _0600_ (.A1(_0065_),
    .A2(_0066_),
    .A3(_0068_),
    .ZN(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _0601_ (.A1(\full_addr[3] ),
    .A2(\full_addr[2] ),
    .Z(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0602_ (.I(_0070_),
    .Z(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _0603_ (.A1(_0048_),
    .A2(_0051_),
    .A3(_0071_),
    .ZN(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__inv_2 _0604_ (.I(\full_addr[3] ),
    .ZN(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _0605_ (.A1(_0073_),
    .A2(_0045_),
    .A3(_0048_),
    .A4(_0050_),
    .ZN(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0606_ (.I(_0074_),
    .Z(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0607_ (.I(_0043_),
    .Z(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0608_ (.I(\full_addr[2] ),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _0609_ (.I(_0077_),
    .Z(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0610_ (.I(_0049_),
    .Z(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _0611_ (.A1(_0076_),
    .A2(_0078_),
    .A3(_0065_),
    .A4(_0079_),
    .ZN(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _0612_ (.A1(_0069_),
    .A2(_0072_),
    .A3(_0075_),
    .A4(_0080_),
    .Z(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0613_ (.A1(_0047_),
    .A2(_0049_),
    .ZN(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0614_ (.A1(_0067_),
    .A2(_0082_),
    .ZN(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0615_ (.I(_0083_),
    .Z(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0616_ (.I(_0084_),
    .Z(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _0617_ (.I(\full_addr[5] ),
    .Z(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _0618_ (.A1(_0055_),
    .A2(_0058_),
    .A3(_0086_),
    .A4(_0060_),
    .ZN(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0619_ (.I(_0087_),
    .Z(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0620_ (.I(_0088_),
    .Z(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_4 _0621_ (.A1(\full_addr[5] ),
    .A2(_0060_),
    .ZN(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _0622_ (.I(\full_addr[7] ),
    .ZN(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0623_ (.I(_0091_),
    .Z(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0624_ (.I(_0037_),
    .Z(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0625_ (.A1(_0092_),
    .A2(_0093_),
    .ZN(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _0626_ (.A1(\full_addr[1] ),
    .A2(\full_addr[0] ),
    .Z(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0627_ (.I(_0095_),
    .Z(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _0628_ (.A1(_0068_),
    .A2(_0096_),
    .Z(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0629_ (.I(_0073_),
    .Z(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0630_ (.I(_0045_),
    .Z(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0631_ (.I(_0064_),
    .Z(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _0632_ (.A1(_0098_),
    .A2(_0099_),
    .A3(_0100_),
    .A4(_0066_),
    .ZN(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0633_ (.I(_0092_),
    .Z(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0634_ (.I(_0059_),
    .Z(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _0635_ (.A1(_0102_),
    .A2(_0093_),
    .A3(_0103_),
    .A4(_0061_),
    .ZN(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _0636_ (.A1(_0090_),
    .A2(_0094_),
    .A3(_0097_),
    .B1(_0101_),
    .B2(_0104_),
    .ZN(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _0637_ (.A1(_0063_),
    .A2(_0081_),
    .B1(_0085_),
    .B2(_0089_),
    .C(_0105_),
    .ZN(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0638_ (.I(_0074_),
    .Z(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _0639_ (.I(_0037_),
    .Z(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _0640_ (.I(\full_addr[4] ),
    .ZN(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _0641_ (.I(_0109_),
    .Z(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _0642_ (.A1(_0036_),
    .A2(_0108_),
    .A3(_0086_),
    .A4(_0110_),
    .ZN(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0643_ (.I(_0111_),
    .Z(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0644_ (.A1(_0107_),
    .A2(_0112_),
    .ZN(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0645_ (.I(_0080_),
    .Z(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _0646_ (.A1(_0055_),
    .A2(_0057_),
    .A3(_0039_),
    .A4(_0109_),
    .ZN(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0647_ (.I(_0115_),
    .Z(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _0648_ (.A1(_0091_),
    .A2(_0108_),
    .A3(_0059_),
    .A4(_0041_),
    .ZN(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _0649_ (.I(_0117_),
    .Z(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0650_ (.I(_0095_),
    .Z(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _0651_ (.A1(_0076_),
    .A2(_0078_),
    .A3(_0119_),
    .ZN(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0652_ (.I(_0120_),
    .Z(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _0653_ (.A1(_0114_),
    .A2(_0116_),
    .B1(_0118_),
    .B2(_0121_),
    .ZN(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _0654_ (.A1(_0091_),
    .A2(_0108_),
    .A3(_0039_),
    .A4(_0060_),
    .ZN(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0655_ (.I(_0123_),
    .Z(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _0656_ (.A1(_0055_),
    .A2(_0108_),
    .A3(_0090_),
    .ZN(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0657_ (.I(_0125_),
    .Z(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _0658_ (.A1(_0068_),
    .A2(_0119_),
    .ZN(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0659_ (.A1(_0124_),
    .A2(_0126_),
    .B(_0127_),
    .ZN(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _0660_ (.A1(_0065_),
    .A2(_0079_),
    .A3(_0071_),
    .ZN(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0661_ (.I(_0129_),
    .Z(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _0662_ (.A1(_0076_),
    .A2(_0077_),
    .A3(_0082_),
    .ZN(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0663_ (.I(_0131_),
    .Z(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0664_ (.I(_0062_),
    .Z(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0665_ (.A1(_0130_),
    .A2(_0132_),
    .B(_0133_),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _0666_ (.A1(_0113_),
    .A2(_0122_),
    .A3(_0128_),
    .A4(_0134_),
    .Z(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _0667_ (.A1(_0048_),
    .A2(_0051_),
    .A3(_0068_),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0668_ (.I(_0136_),
    .Z(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0669_ (.A1(_0124_),
    .A2(_0137_),
    .ZN(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _0670_ (.I(_0083_),
    .Z(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _0671_ (.A1(_0073_),
    .A2(_0046_),
    .A3(_0065_),
    .A4(_0079_),
    .ZN(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0672_ (.I(_0140_),
    .Z(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _0673_ (.A1(_0056_),
    .A2(_0058_),
    .A3(_0090_),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0674_ (.I(_0142_),
    .Z(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _0675_ (.A1(_0139_),
    .A2(_0141_),
    .B(_0143_),
    .ZN(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0676_ (.I(_0123_),
    .Z(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0677_ (.I(_0145_),
    .Z(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0678_ (.I(_0140_),
    .Z(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0679_ (.A1(_0146_),
    .A2(_0147_),
    .ZN(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0680_ (.I(_0142_),
    .Z(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0681_ (.A1(_0107_),
    .A2(_0149_),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _0682_ (.A1(_0138_),
    .A2(_0144_),
    .A3(_0148_),
    .A4(_0150_),
    .Z(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_4 _0683_ (.A1(_0106_),
    .A2(_0135_),
    .A3(_0151_),
    .ZN(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _0684_ (.I(_0140_),
    .Z(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _0685_ (.A1(_0036_),
    .A2(_0038_),
    .A3(_0059_),
    .A4(_0041_),
    .ZN(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0686_ (.I(_0154_),
    .Z(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0687_ (.I(_0076_),
    .Z(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0688_ (.I(_0077_),
    .Z(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0689_ (.I(_0047_),
    .Z(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _0690_ (.A1(_0044_),
    .A2(_0099_),
    .A3(_0158_),
    .A4(_0066_),
    .ZN(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _0691_ (.A1(_0156_),
    .A2(_0157_),
    .A3(_0096_),
    .B(_0159_),
    .ZN(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _0692_ (.A1(_0153_),
    .A2(_0155_),
    .B1(_0160_),
    .B2(_0112_),
    .ZN(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _0693_ (.A1(_0035_),
    .A2(_0042_),
    .A3(_0159_),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0694_ (.A1(\writable[8] ),
    .A2(_0162_),
    .ZN(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _0695_ (.A1(_0043_),
    .A2(_0077_),
    .A3(_0047_),
    .A4(_0050_),
    .ZN(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0696_ (.I(_0164_),
    .Z(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _0697_ (.A1(_0092_),
    .A2(_0038_),
    .A3(_0086_),
    .A4(_0110_),
    .ZN(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _0698_ (.I(_0166_),
    .Z(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _0699_ (.A1(_0165_),
    .A2(_0084_),
    .A3(_0120_),
    .B(_0167_),
    .ZN(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _0700_ (.A1(_0161_),
    .A2(_0163_),
    .A3(_0168_),
    .ZN(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _0701_ (.A1(_0035_),
    .A2(_0042_),
    .A3(_0052_),
    .Z(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0702_ (.I(_0170_),
    .Z(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _0703_ (.A1(_0092_),
    .A2(_0093_),
    .A3(_0090_),
    .ZN(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0704_ (.I(_0172_),
    .Z(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0705_ (.I(_0082_),
    .Z(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _0706_ (.A1(_0119_),
    .A2(_0174_),
    .B(_0098_),
    .C(_0099_),
    .ZN(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0707_ (.I(_0046_),
    .Z(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__or4_2 _0708_ (.A1(\full_addr[7] ),
    .A2(_0037_),
    .A3(\full_addr[5] ),
    .A4(\full_addr[4] ),
    .Z(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0709_ (.I(_0177_),
    .Z(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _0710_ (.A1(_0098_),
    .A2(_0176_),
    .A3(_0096_),
    .A4(_0178_),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0711_ (.I(_0179_),
    .Z(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0712_ (.A1(_0173_),
    .A2(_0175_),
    .B1(_0180_),
    .B2(net15),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0713_ (.I(_0069_),
    .Z(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0714_ (.I(_0117_),
    .Z(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0715_ (.A1(_0071_),
    .A2(_0095_),
    .ZN(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0716_ (.I(_0184_),
    .Z(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0717_ (.I(_0185_),
    .Z(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0718_ (.A1(_0182_),
    .A2(_0183_),
    .B1(_0186_),
    .B2(_0149_),
    .ZN(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _0719_ (.A1(_0171_),
    .A2(_0181_),
    .A3(_0187_),
    .Z(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _0720_ (.I(net12),
    .ZN(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0721_ (.I(_0080_),
    .Z(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _0722_ (.A1(_0036_),
    .A2(_0038_),
    .A3(_0086_),
    .A4(_0041_),
    .ZN(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0723_ (.I(_0191_),
    .Z(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0724_ (.I(_0192_),
    .Z(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0725_ (.A1(net10),
    .A2(net11),
    .ZN(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _0726_ (.A1(_0189_),
    .A2(_0190_),
    .A3(_0193_),
    .A4(_0194_),
    .ZN(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0727_ (.I(_0115_),
    .Z(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0728_ (.I(_0196_),
    .Z(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0729_ (.A1(_0197_),
    .A2(_0085_),
    .ZN(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0730_ (.I(_0072_),
    .Z(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0731_ (.I(_0111_),
    .Z(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0732_ (.I(_0120_),
    .Z(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _0733_ (.A1(_0199_),
    .A2(_0200_),
    .B1(_0201_),
    .B2(_0063_),
    .ZN(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _0734_ (.A1(_0188_),
    .A2(_0195_),
    .A3(_0198_),
    .A4(_0202_),
    .ZN(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0735_ (.A1(_0101_),
    .A2(_0178_),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0736_ (.I(_0204_),
    .Z(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _0737_ (.A1(_0044_),
    .A2(_0078_),
    .A3(_0096_),
    .A4(_0177_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0738_ (.I(_0206_),
    .Z(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0739_ (.I(_0093_),
    .Z(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _0740_ (.A1(_0102_),
    .A2(_0208_),
    .A3(_0040_),
    .A4(_0110_),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0741_ (.A1(_0156_),
    .A2(_0157_),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _0742_ (.A1(_0056_),
    .A2(_0058_),
    .A3(_0040_),
    .A4(_0110_),
    .ZN(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_4 _0743_ (.A1(_0209_),
    .A2(_0210_),
    .A3(_0174_),
    .B1(_0211_),
    .B2(_0097_),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _0744_ (.A1(net31),
    .A2(_0205_),
    .B1(_0207_),
    .B2(net45),
    .C(_0212_),
    .ZN(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0745_ (.A1(_0072_),
    .A2(_0087_),
    .ZN(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0746_ (.I(_0165_),
    .Z(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0747_ (.A1(_0215_),
    .A2(_0089_),
    .ZN(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _0748_ (.A1(_0044_),
    .A2(_0078_),
    .A3(_0174_),
    .A4(_0178_),
    .ZN(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0749_ (.I(_0217_),
    .Z(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0750_ (.A1(net29),
    .A2(_0218_),
    .ZN(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _0751_ (.A1(_0214_),
    .A2(_0216_),
    .A3(_0219_),
    .Z(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0752_ (.I(_0136_),
    .Z(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0753_ (.A1(_0073_),
    .A2(_0046_),
    .A3(_0119_),
    .ZN(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0754_ (.I(_0222_),
    .Z(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0755_ (.I(_0223_),
    .Z(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_4 _0756_ (.A1(_0221_),
    .A2(_0224_),
    .B(_0063_),
    .ZN(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _0757_ (.I(_0196_),
    .Z(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0758_ (.I(_0153_),
    .Z(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0759_ (.I(_0191_),
    .Z(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _0760_ (.A1(_0182_),
    .A2(_0226_),
    .B1(_0227_),
    .B2(_0228_),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _0761_ (.A1(_0213_),
    .A2(_0220_),
    .A3(_0225_),
    .A4(_0229_),
    .ZN(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _0762_ (.A1(_0152_),
    .A2(_0169_),
    .A3(_0203_),
    .A4(_0230_),
    .ZN(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0763_ (.I(_0127_),
    .Z(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0764_ (.A1(_0116_),
    .A2(_0232_),
    .ZN(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _0765_ (.A1(_0127_),
    .A2(_0112_),
    .B1(_0185_),
    .B2(_0088_),
    .C1(_0153_),
    .C2(_0196_),
    .ZN(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _0766_ (.I(_0129_),
    .Z(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0767_ (.I(_0222_),
    .Z(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0768_ (.I(_0125_),
    .Z(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0769_ (.A1(_0235_),
    .A2(_0236_),
    .B(_0237_),
    .ZN(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0770_ (.I(_0131_),
    .Z(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0771_ (.A1(_0121_),
    .A2(_0239_),
    .B(_0154_),
    .ZN(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _0772_ (.A1(_0233_),
    .A2(_0234_),
    .A3(_0238_),
    .A4(_0240_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0773_ (.I(_0120_),
    .Z(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0774_ (.I(_0172_),
    .Z(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0775_ (.A1(_0242_),
    .A2(_0243_),
    .ZN(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0776_ (.I(_0164_),
    .Z(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _0777_ (.A1(_0114_),
    .A2(_0167_),
    .B1(_0243_),
    .B2(_0245_),
    .ZN(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0778_ (.I(_0184_),
    .Z(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _0779_ (.A1(_0121_),
    .A2(_0237_),
    .B1(_0243_),
    .B2(_0247_),
    .C1(_0154_),
    .C2(_0139_),
    .ZN(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0780_ (.A1(_0098_),
    .A2(_0099_),
    .A3(_0174_),
    .ZN(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0781_ (.I(_0249_),
    .Z(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _0782_ (.A1(_0102_),
    .A2(_0208_),
    .A3(_0103_),
    .ZN(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _0783_ (.A1(_0118_),
    .A2(_0223_),
    .B1(_0250_),
    .B2(_0167_),
    .C1(_0251_),
    .C2(_0114_),
    .ZN(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _0784_ (.A1(_0244_),
    .A2(_0246_),
    .A3(_0248_),
    .A4(_0252_),
    .ZN(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0785_ (.I(_0249_),
    .Z(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0786_ (.A1(_0146_),
    .A2(_0126_),
    .B(_0254_),
    .ZN(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0787_ (.I(_0117_),
    .Z(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _0788_ (.A1(_0143_),
    .A2(_0130_),
    .B1(_0239_),
    .B2(_0256_),
    .C1(_0167_),
    .C2(_0127_),
    .ZN(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0789_ (.A1(_0255_),
    .A2(_0257_),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0790_ (.I(_0069_),
    .Z(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0791_ (.I(_0166_),
    .Z(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0792_ (.A1(_0259_),
    .A2(_0199_),
    .B(_0260_),
    .ZN(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _0793_ (.A1(_0075_),
    .A2(_0118_),
    .B1(_0235_),
    .B2(_0192_),
    .C1(_0250_),
    .C2(_0142_),
    .ZN(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0794_ (.A1(_0261_),
    .A2(_0262_),
    .ZN(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _0795_ (.A1(_0241_),
    .A2(_0253_),
    .A3(_0258_),
    .A4(_0263_),
    .ZN(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0796_ (.A1(_0070_),
    .A2(_0082_),
    .ZN(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0797_ (.I(_0265_),
    .Z(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0798_ (.I(_0266_),
    .Z(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0799_ (.A1(_0197_),
    .A2(_0193_),
    .B(_0267_),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0800_ (.I(_0087_),
    .Z(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0801_ (.A1(_0075_),
    .A2(_0269_),
    .ZN(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _0802_ (.A1(_0165_),
    .A2(_0175_),
    .A3(_0185_),
    .B(_0154_),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _0803_ (.A1(_0157_),
    .A2(_0100_),
    .A3(_0066_),
    .ZN(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0804_ (.A1(_0185_),
    .A2(_0272_),
    .B(_0237_),
    .ZN(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0805_ (.A1(_0196_),
    .A2(_0223_),
    .ZN(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _0806_ (.A1(_0157_),
    .A2(_0158_),
    .A3(_0051_),
    .ZN(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0807_ (.I(_0079_),
    .Z(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _0808_ (.A1(_0176_),
    .A2(_0100_),
    .A3(_0276_),
    .ZN(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0809_ (.A1(_0275_),
    .A2(_0277_),
    .B(_0112_),
    .ZN(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__and4_2 _0810_ (.A1(_0271_),
    .A2(_0273_),
    .A3(_0274_),
    .A4(_0278_),
    .Z(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0811_ (.I(_0279_),
    .Z(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _0812_ (.A1(_0264_),
    .A2(_0268_),
    .A3(_0270_),
    .A4(_0280_),
    .Z(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _0813_ (.A1(_0032_),
    .A2(_0054_),
    .B1(_0231_),
    .B2(_0281_),
    .ZN(net49));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0814_ (.I(\writable[1] ),
    .ZN(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0815_ (.A1(_0106_),
    .A2(_0135_),
    .ZN(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0816_ (.A1(_0270_),
    .A2(_0280_),
    .ZN(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0817_ (.I(\writable[9] ),
    .ZN(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _0818_ (.A1(_0035_),
    .A2(_0042_),
    .A3(_0159_),
    .Z(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0819_ (.A1(_0139_),
    .A2(_0141_),
    .B(_0133_),
    .ZN(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0820_ (.A1(_0136_),
    .A2(_0247_),
    .B(_0116_),
    .ZN(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _0821_ (.A1(_0285_),
    .A2(_0286_),
    .B(_0287_),
    .C(_0288_),
    .ZN(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _0822_ (.A1(_0189_),
    .A2(_0190_),
    .A3(_0192_),
    .ZN(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0823_ (.I(net11),
    .ZN(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0824_ (.A1(net10),
    .A2(_0291_),
    .ZN(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0825_ (.I(_0166_),
    .Z(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _0826_ (.A1(_0259_),
    .A2(_0256_),
    .B1(_0242_),
    .B2(_0293_),
    .ZN(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _0827_ (.A1(_0084_),
    .A2(_0145_),
    .B1(_0125_),
    .B2(_0074_),
    .ZN(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _0828_ (.A1(_0290_),
    .A2(_0292_),
    .B(_0294_),
    .C(_0295_),
    .ZN(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0829_ (.I(_0206_),
    .Z(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0830_ (.A1(net46),
    .A2(_0297_),
    .B1(_0218_),
    .B2(net30),
    .ZN(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0831_ (.A1(net22),
    .A2(_0180_),
    .ZN(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0832_ (.A1(_0171_),
    .A2(_0298_),
    .A3(_0299_),
    .ZN(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _0833_ (.A1(_0143_),
    .A2(_0242_),
    .B1(_0137_),
    .B2(_0293_),
    .C1(_0247_),
    .C2(_0124_),
    .ZN(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0834_ (.I(_0191_),
    .Z(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0835_ (.A1(_0139_),
    .A2(_0260_),
    .B1(_0302_),
    .B2(_0147_),
    .ZN(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0836_ (.A1(_0107_),
    .A2(_0173_),
    .ZN(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0837_ (.I(_0145_),
    .Z(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0838_ (.A1(_0190_),
    .A2(_0305_),
    .ZN(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _0839_ (.A1(_0301_),
    .A2(_0303_),
    .A3(_0304_),
    .A4(_0306_),
    .ZN(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _0840_ (.A1(_0289_),
    .A2(_0296_),
    .A3(_0300_),
    .A4(_0307_),
    .Z(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0841_ (.A1(_0103_),
    .A2(_0061_),
    .ZN(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0842_ (.A1(_0103_),
    .A2(_0075_),
    .B1(_0130_),
    .B2(_0309_),
    .ZN(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0843_ (.A1(_0126_),
    .A2(_0266_),
    .ZN(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _0844_ (.A1(_0102_),
    .A2(_0208_),
    .A3(_0310_),
    .B(_0311_),
    .ZN(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _0845_ (.A1(_0156_),
    .A2(_0176_),
    .A3(_0100_),
    .A4(_0276_),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0846_ (.A1(_0313_),
    .A2(_0178_),
    .B(_0161_),
    .ZN(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _0847_ (.A1(_0293_),
    .A2(_0247_),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _0848_ (.A1(_0237_),
    .A2(_0153_),
    .B1(_0172_),
    .B2(_0235_),
    .ZN(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _0849_ (.A1(_0138_),
    .A2(_0144_),
    .A3(_0315_),
    .A4(_0316_),
    .ZN(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0850_ (.A1(net38),
    .A2(_0245_),
    .A3(_0302_),
    .ZN(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0851_ (.A1(_0269_),
    .A2(_0266_),
    .ZN(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0852_ (.A1(_0084_),
    .A2(_0191_),
    .B1(_0265_),
    .B2(_0145_),
    .ZN(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0853_ (.I(_0320_),
    .Z(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _0854_ (.A1(_0214_),
    .A2(_0318_),
    .A3(_0319_),
    .A4(_0321_),
    .ZN(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _0855_ (.A1(_0312_),
    .A2(_0314_),
    .A3(_0317_),
    .A4(_0322_),
    .Z(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _0856_ (.A1(_0283_),
    .A2(_0284_),
    .A3(_0308_),
    .A4(_0323_),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _0857_ (.A1(_0282_),
    .A2(_0054_),
    .B1(_0264_),
    .B2(_0324_),
    .ZN(net50));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0858_ (.I(\writable[2] ),
    .ZN(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0859_ (.A1(_0245_),
    .A2(_0186_),
    .B(_0143_),
    .ZN(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _0860_ (.A1(_0287_),
    .A2(_0288_),
    .A3(_0326_),
    .ZN(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0861_ (.A1(_0245_),
    .A2(_0254_),
    .B(_0256_),
    .ZN(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0862_ (.A1(_0141_),
    .A2(_0260_),
    .B1(_0186_),
    .B2(_0200_),
    .ZN(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0863_ (.A1(_0328_),
    .A2(_0329_),
    .ZN(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0864_ (.A1(_0212_),
    .A2(_0327_),
    .A3(_0330_),
    .ZN(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0865_ (.I(_0179_),
    .Z(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _0866_ (.A1(net23),
    .A2(_0332_),
    .B1(_0205_),
    .B2(net39),
    .C1(_0207_),
    .C2(net32),
    .ZN(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0867_ (.I(_0214_),
    .Z(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0868_ (.A1(_0334_),
    .A2(_0319_),
    .ZN(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0869_ (.A1(_0259_),
    .A2(_0116_),
    .ZN(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _0870_ (.A1(_0124_),
    .A2(_0239_),
    .B1(_0223_),
    .B2(_0088_),
    .ZN(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0871_ (.A1(net16),
    .A2(_0218_),
    .ZN(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0872_ (.I(_0266_),
    .Z(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0873_ (.A1(_0133_),
    .A2(_0339_),
    .ZN(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _0874_ (.A1(_0336_),
    .A2(_0337_),
    .A3(_0338_),
    .A4(_0340_),
    .ZN(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _0875_ (.A1(_0183_),
    .A2(_0137_),
    .B1(_0173_),
    .B2(_0339_),
    .ZN(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0876_ (.I(_0118_),
    .Z(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0877_ (.A1(_0085_),
    .A2(_0343_),
    .ZN(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0878_ (.I(_0235_),
    .Z(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0879_ (.I(_0166_),
    .Z(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0880_ (.A1(_0215_),
    .A2(_0345_),
    .B(_0346_),
    .ZN(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0881_ (.I(_0142_),
    .Z(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0882_ (.I(_0074_),
    .Z(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0883_ (.A1(_0226_),
    .A2(_0232_),
    .B1(_0348_),
    .B2(_0349_),
    .ZN(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _0884_ (.A1(_0342_),
    .A2(_0344_),
    .A3(_0347_),
    .A4(_0350_),
    .ZN(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _0885_ (.A1(_0258_),
    .A2(_0335_),
    .A3(_0341_),
    .A4(_0351_),
    .ZN(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0886_ (.A1(_0158_),
    .A2(_0071_),
    .ZN(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0887_ (.A1(_0305_),
    .A2(_0353_),
    .ZN(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0888_ (.A1(_0321_),
    .A2(_0354_),
    .ZN(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0889_ (.I(net10),
    .Z(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0890_ (.A1(_0356_),
    .A2(_0291_),
    .A3(_0290_),
    .ZN(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0891_ (.A1(_0161_),
    .A2(_0244_),
    .A3(_0246_),
    .ZN(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0892_ (.A1(_0355_),
    .A2(_0357_),
    .A3(_0358_),
    .ZN(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _0893_ (.A1(_0331_),
    .A2(_0333_),
    .A3(_0352_),
    .A4(_0359_),
    .Z(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _0894_ (.A1(_0268_),
    .A2(_0270_),
    .A3(_0280_),
    .ZN(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _0895_ (.A1(_0113_),
    .A2(_0122_),
    .A3(_0128_),
    .A4(_0134_),
    .ZN(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0896_ (.A1(_0343_),
    .A2(_0267_),
    .Z(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0897_ (.A1(_0269_),
    .A2(_0254_),
    .ZN(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _0898_ (.A1(_0199_),
    .A2(_0226_),
    .B1(_0132_),
    .B2(_0293_),
    .ZN(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0899_ (.A1(_0133_),
    .A2(_0183_),
    .B(_0186_),
    .ZN(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _0900_ (.A1(_0364_),
    .A2(_0365_),
    .A3(_0366_),
    .ZN(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _0901_ (.A1(_0362_),
    .A2(_0312_),
    .A3(_0363_),
    .A4(_0367_),
    .Z(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0902_ (.I(_0165_),
    .Z(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _0903_ (.A1(_0121_),
    .A2(_0250_),
    .Z(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _0904_ (.I(_0088_),
    .Z(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_4 _0905_ (.A1(_0063_),
    .A2(_0369_),
    .B1(_0370_),
    .B2(_0226_),
    .C1(_0371_),
    .C2(_0182_),
    .ZN(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _0906_ (.A1(_0149_),
    .A2(_0146_),
    .A3(_0155_),
    .B(_0259_),
    .ZN(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0907_ (.A1(_0200_),
    .A2(_0236_),
    .B1(_0339_),
    .B2(_0155_),
    .ZN(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0908_ (.A1(_0089_),
    .A2(_0137_),
    .B1(_0254_),
    .B2(_0302_),
    .ZN(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _0909_ (.A1(_0373_),
    .A2(_0374_),
    .A3(_0375_),
    .Z(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _0910_ (.A1(_0106_),
    .A2(_0225_),
    .A3(_0372_),
    .A4(_0376_),
    .ZN(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0911_ (.I(_0170_),
    .Z(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0912_ (.I(_0162_),
    .Z(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0913_ (.A1(\writable[10] ),
    .A2(_0379_),
    .ZN(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0914_ (.A1(_0378_),
    .A2(_0380_),
    .ZN(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _0915_ (.A1(_0361_),
    .A2(_0368_),
    .A3(_0377_),
    .A4(_0381_),
    .ZN(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _0916_ (.A1(_0325_),
    .A2(_0054_),
    .B1(_0360_),
    .B2(_0382_),
    .ZN(net51));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0917_ (.I(\writable[3] ),
    .ZN(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0918_ (.I(_0280_),
    .ZN(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0919_ (.A1(_0225_),
    .A2(_0372_),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _0920_ (.A1(_0241_),
    .A2(_0384_),
    .A3(_0367_),
    .A4(_0385_),
    .ZN(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0921_ (.A1(_0106_),
    .A2(_0135_),
    .Z(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0922_ (.A1(_0224_),
    .A2(_0267_),
    .B(_0149_),
    .ZN(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0923_ (.A1(_0215_),
    .A2(_0305_),
    .B1(_0173_),
    .B2(_0199_),
    .ZN(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0924_ (.A1(_0201_),
    .A2(_0132_),
    .B(_0269_),
    .ZN(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0925_ (.A1(_0388_),
    .A2(_0389_),
    .A3(_0390_),
    .ZN(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _0926_ (.A1(_0263_),
    .A2(_0327_),
    .A3(_0391_),
    .ZN(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _0927_ (.A1(_0138_),
    .A2(_0144_),
    .A3(_0148_),
    .ZN(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0928_ (.A1(_0256_),
    .A2(_0141_),
    .ZN(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0929_ (.A1(_0089_),
    .A2(_0147_),
    .B1(_0228_),
    .B2(_0182_),
    .ZN(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0930_ (.A1(_0221_),
    .A2(_0346_),
    .B1(_0224_),
    .B2(_0343_),
    .ZN(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _0931_ (.A1(_0378_),
    .A2(_0394_),
    .A3(_0395_),
    .A4(_0396_),
    .ZN(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0932_ (.A1(_0369_),
    .A2(_0201_),
    .B(_0346_),
    .ZN(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _0933_ (.A1(net24),
    .A2(_0180_),
    .B1(_0297_),
    .B2(net33),
    .ZN(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _0934_ (.A1(_0398_),
    .A2(_0334_),
    .A3(_0216_),
    .A4(_0399_),
    .ZN(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _0935_ (.I(_0217_),
    .Z(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0936_ (.A1(net17),
    .A2(_0401_),
    .ZN(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0937_ (.I(_0239_),
    .Z(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _0938_ (.I(_0172_),
    .Z(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0939_ (.A1(_0403_),
    .A2(_0224_),
    .B(_0404_),
    .ZN(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0940_ (.A1(_0349_),
    .A2(_0403_),
    .B(_0348_),
    .ZN(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0941_ (.A1(net40),
    .A2(_0369_),
    .A3(_0228_),
    .ZN(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _0942_ (.A1(_0402_),
    .A2(_0405_),
    .A3(_0406_),
    .A4(_0407_),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _0943_ (.A1(_0393_),
    .A2(_0397_),
    .A3(_0400_),
    .A4(_0408_),
    .ZN(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _0944_ (.I(_0295_),
    .Z(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0945_ (.A1(_0345_),
    .A2(_0346_),
    .ZN(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _0946_ (.A1(_0410_),
    .A2(_0315_),
    .A3(_0316_),
    .A4(_0411_),
    .ZN(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0947_ (.A1(net10),
    .A2(net11),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0948_ (.A1(_0290_),
    .A2(_0413_),
    .ZN(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _0949_ (.A1(\writable[11] ),
    .A2(_0379_),
    .B(_0412_),
    .C(_0414_),
    .ZN(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _0950_ (.A1(_0387_),
    .A2(_0392_),
    .A3(_0409_),
    .A4(_0415_),
    .Z(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _0951_ (.A1(_0383_),
    .A2(_0054_),
    .B1(_0386_),
    .B2(_0416_),
    .ZN(net52));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _0952_ (.I(\writable[4] ),
    .ZN(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__buf_3 _0953_ (.I(_0053_),
    .Z(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _0954_ (.A1(net12),
    .A2(_0114_),
    .A3(_0192_),
    .Z(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _0955_ (.A1(_0287_),
    .A2(_0288_),
    .A3(_0321_),
    .A4(_0354_),
    .ZN(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _0956_ (.A1(\writable[12] ),
    .A2(_0379_),
    .B1(_0194_),
    .B2(_0419_),
    .C(_0420_),
    .ZN(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0957_ (.A1(_0215_),
    .A2(_0267_),
    .B(_0371_),
    .ZN(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _0958_ (.A1(_0246_),
    .A2(_0410_),
    .A3(_0337_),
    .A4(_0422_),
    .ZN(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0959_ (.A1(_0197_),
    .A2(_0232_),
    .B1(_0227_),
    .B2(_0404_),
    .ZN(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _0960_ (.A1(_0378_),
    .A2(_0229_),
    .A3(_0304_),
    .A4(_0424_),
    .ZN(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0961_ (.A1(net41),
    .A2(_0369_),
    .A3(_0193_),
    .ZN(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0962_ (.A1(net18),
    .A2(_0401_),
    .ZN(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _0963_ (.A1(net25),
    .A2(_0332_),
    .B1(_0297_),
    .B2(net34),
    .ZN(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0964_ (.A1(_0426_),
    .A2(_0427_),
    .A3(_0428_),
    .ZN(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _0965_ (.A1(_0263_),
    .A2(_0423_),
    .A3(_0425_),
    .A4(_0429_),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _0966_ (.A1(_0421_),
    .A2(_0430_),
    .Z(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _0967_ (.A1(_0168_),
    .A2(_0328_),
    .A3(_0329_),
    .Z(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _0968_ (.A1(_0315_),
    .A2(_0316_),
    .A3(_0342_),
    .A4(_0432_),
    .ZN(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _0969_ (.A1(_0314_),
    .A2(_0391_),
    .Z(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _0970_ (.A1(_0152_),
    .A2(_0284_),
    .A3(_0433_),
    .A4(_0434_),
    .ZN(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _0971_ (.A1(_0417_),
    .A2(_0418_),
    .B1(_0431_),
    .B2(_0435_),
    .ZN(net53));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _0972_ (.I(\writable[5] ),
    .ZN(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _0973_ (.A1(_0362_),
    .A2(_0363_),
    .ZN(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _0974_ (.A1(_0348_),
    .A2(_0201_),
    .B(_0327_),
    .ZN(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0975_ (.A1(_0356_),
    .A2(_0291_),
    .A3(_0419_),
    .ZN(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0976_ (.A1(_0243_),
    .A2(_0250_),
    .ZN(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _0977_ (.A1(_0168_),
    .A2(_0336_),
    .A3(_0320_),
    .A4(_0440_),
    .Z(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _0978_ (.A1(_0410_),
    .A2(_0411_),
    .A3(_0439_),
    .A4(_0441_),
    .Z(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _0979_ (.A1(_0276_),
    .A2(_0146_),
    .A3(_0353_),
    .ZN(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _0980_ (.A1(_0349_),
    .A2(_0371_),
    .B1(_0343_),
    .B2(_0227_),
    .C1(_0180_),
    .C2(net26),
    .ZN(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _0981_ (.A1(net42),
    .A2(_0204_),
    .B1(_0297_),
    .B2(net35),
    .C1(_0218_),
    .C2(net19),
    .ZN(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _0982_ (.A1(_0337_),
    .A2(_0443_),
    .A3(_0444_),
    .A4(_0445_),
    .Z(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _0983_ (.A1(_0437_),
    .A2(_0438_),
    .A3(_0442_),
    .A4(_0446_),
    .Z(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _0984_ (.A1(_0234_),
    .A2(_0238_),
    .A3(_0240_),
    .Z(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _0985_ (.A1(_0345_),
    .A2(_0221_),
    .B(_0155_),
    .ZN(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0986_ (.A1(_0200_),
    .A2(_0403_),
    .ZN(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _0987_ (.A1(_0334_),
    .A2(_0449_),
    .A3(_0450_),
    .Z(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _0988_ (.A1(_0448_),
    .A2(_0422_),
    .A3(_0451_),
    .ZN(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _0989_ (.A1(_0349_),
    .A2(_0232_),
    .B(_0193_),
    .ZN(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0990_ (.A1(_0371_),
    .A2(_0345_),
    .ZN(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _0991_ (.A1(_0197_),
    .A2(_0403_),
    .B1(_0275_),
    .B2(_0126_),
    .ZN(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _0992_ (.A1(_0279_),
    .A2(_0453_),
    .A3(_0454_),
    .A4(_0455_),
    .ZN(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0993_ (.A1(\writable[13] ),
    .A2(_0379_),
    .ZN(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _0994_ (.A1(_0378_),
    .A2(_0457_),
    .ZN(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _0995_ (.A1(_0317_),
    .A2(_0452_),
    .A3(_0456_),
    .A4(_0458_),
    .ZN(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _0996_ (.A1(_0436_),
    .A2(_0418_),
    .B1(_0447_),
    .B2(_0459_),
    .ZN(net54));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _0997_ (.I(\writable[6] ),
    .ZN(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _0998_ (.A1(_0209_),
    .A2(_0313_),
    .B(_0372_),
    .C(_0135_),
    .ZN(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _0999_ (.A1(_0433_),
    .A2(_0461_),
    .ZN(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1000_ (.A1(_0410_),
    .A2(_0321_),
    .ZN(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1001_ (.A1(_0334_),
    .A2(_0336_),
    .ZN(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _1002_ (.A1(_0242_),
    .A2(_0130_),
    .A3(_0236_),
    .B(_0305_),
    .ZN(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1003_ (.A1(_0085_),
    .A2(_0183_),
    .B1(_0147_),
    .B2(_0404_),
    .ZN(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1004_ (.A1(_0150_),
    .A2(_0411_),
    .A3(_0465_),
    .A4(_0466_),
    .ZN(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _1005_ (.A1(_0053_),
    .A2(_0463_),
    .A3(_0464_),
    .A4(_0467_),
    .ZN(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _1006_ (.A1(_0260_),
    .A2(_0339_),
    .B1(_0353_),
    .B2(_0302_),
    .ZN(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1007_ (.A1(net27),
    .A2(_0332_),
    .B1(_0401_),
    .B2(net20),
    .ZN(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1008_ (.A1(net43),
    .A2(_0205_),
    .B1(_0207_),
    .B2(net36),
    .ZN(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _1009_ (.A1(_0270_),
    .A2(_0337_),
    .A3(_0394_),
    .Z(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1010_ (.A1(_0469_),
    .A2(_0470_),
    .A3(_0471_),
    .A4(_0472_),
    .Z(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1011_ (.A1(_0356_),
    .A2(_0291_),
    .ZN(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _1012_ (.A1(_0107_),
    .A2(_0190_),
    .A3(_0132_),
    .A4(_0236_),
    .Z(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _1013_ (.A1(\writable[14] ),
    .A2(_0162_),
    .B1(_0474_),
    .B2(_0419_),
    .C1(_0475_),
    .C2(_0404_),
    .ZN(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _1014_ (.A1(_0438_),
    .A2(_0468_),
    .A3(_0473_),
    .A4(_0476_),
    .Z(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _1015_ (.A1(_0460_),
    .A2(_0418_),
    .B1(_0462_),
    .B2(_0477_),
    .ZN(net55));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1016_ (.I(\writable[7] ),
    .ZN(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1017_ (.A1(_0212_),
    .A2(_0327_),
    .A3(_0330_),
    .Z(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _1018_ (.A1(_0479_),
    .A2(_0434_),
    .A3(_0461_),
    .ZN(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1019_ (.A1(_0356_),
    .A2(net11),
    .A3(_0419_),
    .ZN(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1020_ (.A1(\writable[15] ),
    .A2(_0162_),
    .ZN(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _1021_ (.A1(_0451_),
    .A2(_0481_),
    .A3(_0482_),
    .ZN(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1022_ (.A1(_0227_),
    .A2(_0228_),
    .ZN(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1023_ (.A1(_0171_),
    .A2(_0484_),
    .A3(_0244_),
    .ZN(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1024_ (.A1(_0348_),
    .A2(_0221_),
    .ZN(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _1025_ (.A1(_0319_),
    .A2(_0340_),
    .A3(_0486_),
    .ZN(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _1026_ (.A1(_0294_),
    .A2(_0295_),
    .A3(_0443_),
    .A4(_0469_),
    .ZN(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _1027_ (.A1(_0485_),
    .A2(_0487_),
    .A3(_0488_),
    .Z(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1028_ (.A1(net28),
    .A2(_0332_),
    .B1(_0401_),
    .B2(net21),
    .ZN(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _1029_ (.A1(net44),
    .A2(_0205_),
    .B1(_0207_),
    .B2(net37),
    .ZN(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _1030_ (.A1(_0490_),
    .A2(_0491_),
    .ZN(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _1031_ (.A1(_0241_),
    .A2(_0483_),
    .A3(_0489_),
    .A4(_0492_),
    .ZN(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_4 _1032_ (.A1(_0478_),
    .A2(_0418_),
    .B1(_0480_),
    .B2(_0493_),
    .ZN(net56));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1033_ (.I(net2),
    .ZN(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1034_ (.I(net14),
    .Z(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _1035_ (.I(net48),
    .ZN(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _1036_ (.A1(_0496_),
    .A2(net47),
    .ZN(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1037_ (.I(_0497_),
    .Z(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1038_ (.I(net14),
    .Z(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1039_ (.A1(_0499_),
    .A2(_0276_),
    .ZN(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1040_ (.A1(_0494_),
    .A2(_0495_),
    .B(_0498_),
    .C(_0500_),
    .ZN(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1041_ (.I(net3),
    .ZN(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1042_ (.A1(_0499_),
    .A2(_0158_),
    .ZN(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1043_ (.A1(_0501_),
    .A2(_0495_),
    .B(_0498_),
    .C(_0502_),
    .ZN(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1044_ (.I(net4),
    .ZN(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1045_ (.A1(_0499_),
    .A2(_0176_),
    .ZN(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1046_ (.A1(_0503_),
    .A2(_0495_),
    .B(_0498_),
    .C(_0504_),
    .ZN(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _1047_ (.I(net5),
    .ZN(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1048_ (.I(net14),
    .Z(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1049_ (.A1(_0506_),
    .A2(_0156_),
    .ZN(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1050_ (.A1(_0505_),
    .A2(_0495_),
    .B(_0498_),
    .C(_0507_),
    .ZN(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1051_ (.I(net6),
    .ZN(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1052_ (.I(net14),
    .Z(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1053_ (.I(_0497_),
    .Z(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1054_ (.A1(_0506_),
    .A2(_0061_),
    .ZN(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1055_ (.A1(_0508_),
    .A2(_0509_),
    .B(_0510_),
    .C(_0511_),
    .ZN(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1056_ (.I(net7),
    .ZN(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1057_ (.A1(_0506_),
    .A2(_0040_),
    .ZN(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1058_ (.A1(_0512_),
    .A2(_0509_),
    .B(_0510_),
    .C(_0513_),
    .ZN(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1059_ (.I(net8),
    .ZN(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1060_ (.A1(_0506_),
    .A2(_0208_),
    .ZN(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1061_ (.A1(_0514_),
    .A2(_0509_),
    .B(_0510_),
    .C(_0515_),
    .ZN(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _1062_ (.I(net9),
    .ZN(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1063_ (.A1(_0056_),
    .A2(_0499_),
    .ZN(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1064_ (.A1(_0516_),
    .A2(_0509_),
    .B(_0510_),
    .C(_0517_),
    .ZN(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1065_ (.A1(net1),
    .A2(_0171_),
    .ZN(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1066_ (.I(_0518_),
    .Z(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1067_ (.I(_0518_),
    .Z(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1068_ (.I(_0496_),
    .Z(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1069_ (.I(_0521_),
    .Z(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1070_ (.A1(\writable[0] ),
    .A2(_0520_),
    .B(_0522_),
    .ZN(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1071_ (.A1(_0494_),
    .A2(_0519_),
    .B(_0523_),
    .ZN(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1072_ (.A1(\writable[1] ),
    .A2(_0520_),
    .B(_0522_),
    .ZN(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1073_ (.A1(_0501_),
    .A2(_0519_),
    .B(_0524_),
    .ZN(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1074_ (.A1(\writable[2] ),
    .A2(_0520_),
    .B(_0522_),
    .ZN(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1075_ (.A1(_0503_),
    .A2(_0519_),
    .B(_0525_),
    .ZN(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1076_ (.A1(\writable[3] ),
    .A2(_0520_),
    .B(_0522_),
    .ZN(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1077_ (.A1(_0505_),
    .A2(_0519_),
    .B(_0526_),
    .ZN(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1078_ (.I(_0518_),
    .Z(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1079_ (.I(_0518_),
    .Z(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1080_ (.I(_0521_),
    .Z(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1081_ (.A1(\writable[4] ),
    .A2(_0528_),
    .B(_0529_),
    .ZN(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1082_ (.A1(_0508_),
    .A2(_0527_),
    .B(_0530_),
    .ZN(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1083_ (.A1(\writable[5] ),
    .A2(_0528_),
    .B(_0529_),
    .ZN(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1084_ (.A1(_0512_),
    .A2(_0527_),
    .B(_0531_),
    .ZN(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1085_ (.A1(\writable[6] ),
    .A2(_0528_),
    .B(_0529_),
    .ZN(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1086_ (.A1(_0514_),
    .A2(_0527_),
    .B(_0532_),
    .ZN(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1087_ (.A1(\writable[7] ),
    .A2(_0528_),
    .B(_0529_),
    .ZN(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1088_ (.A1(_0516_),
    .A2(_0527_),
    .B(_0533_),
    .ZN(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1089_ (.I(net13),
    .Z(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1090_ (.I(_0497_),
    .Z(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1091_ (.I(net13),
    .Z(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1092_ (.A1(_0536_),
    .A2(\full_addr[8] ),
    .ZN(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1093_ (.A1(_0494_),
    .A2(_0534_),
    .B(_0535_),
    .C(_0537_),
    .ZN(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1094_ (.A1(_0536_),
    .A2(\full_addr[9] ),
    .ZN(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1095_ (.A1(_0501_),
    .A2(_0534_),
    .B(_0535_),
    .C(_0538_),
    .ZN(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1096_ (.A1(_0536_),
    .A2(\full_addr[10] ),
    .ZN(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1097_ (.A1(_0503_),
    .A2(_0534_),
    .B(_0535_),
    .C(_0539_),
    .ZN(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1098_ (.I(net13),
    .Z(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1099_ (.A1(_0540_),
    .A2(\full_addr[11] ),
    .ZN(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1100_ (.A1(_0505_),
    .A2(_0534_),
    .B(_0535_),
    .C(_0541_),
    .ZN(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1101_ (.I(net13),
    .Z(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _1102_ (.I(_0497_),
    .Z(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1103_ (.A1(_0540_),
    .A2(\full_addr[12] ),
    .ZN(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1104_ (.A1(_0508_),
    .A2(_0542_),
    .B(_0543_),
    .C(_0544_),
    .ZN(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1105_ (.A1(_0540_),
    .A2(\full_addr[13] ),
    .ZN(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1106_ (.A1(_0512_),
    .A2(_0542_),
    .B(_0543_),
    .C(_0545_),
    .ZN(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1107_ (.A1(_0540_),
    .A2(\full_addr[14] ),
    .ZN(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1108_ (.A1(_0514_),
    .A2(_0542_),
    .B(_0543_),
    .C(_0546_),
    .ZN(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _1109_ (.A1(\full_addr[15] ),
    .A2(_0536_),
    .ZN(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _1110_ (.A1(_0516_),
    .A2(_0542_),
    .B(_0543_),
    .C(_0547_),
    .ZN(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _1111_ (.A1(net1),
    .A2(_0286_),
    .ZN(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1112_ (.I(_0548_),
    .Z(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1113_ (.I(_0548_),
    .Z(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1114_ (.I(_0521_),
    .Z(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1115_ (.A1(\writable[8] ),
    .A2(_0550_),
    .B(_0551_),
    .ZN(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1116_ (.A1(_0494_),
    .A2(_0549_),
    .B(_0552_),
    .ZN(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1117_ (.A1(\writable[9] ),
    .A2(_0550_),
    .B(_0551_),
    .ZN(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1118_ (.A1(_0501_),
    .A2(_0549_),
    .B(_0553_),
    .ZN(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1119_ (.A1(\writable[10] ),
    .A2(_0550_),
    .B(_0551_),
    .ZN(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1120_ (.A1(_0503_),
    .A2(_0549_),
    .B(_0554_),
    .ZN(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1121_ (.A1(\writable[11] ),
    .A2(_0550_),
    .B(_0551_),
    .ZN(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1122_ (.A1(_0505_),
    .A2(_0549_),
    .B(_0555_),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1123_ (.I(_0548_),
    .Z(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1124_ (.I(_0548_),
    .Z(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _1125_ (.I(_0521_),
    .Z(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1126_ (.A1(\writable[12] ),
    .A2(_0557_),
    .B(_0558_),
    .ZN(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1127_ (.A1(_0508_),
    .A2(_0556_),
    .B(_0559_),
    .ZN(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1128_ (.A1(\writable[13] ),
    .A2(_0557_),
    .B(_0558_),
    .ZN(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1129_ (.A1(_0512_),
    .A2(_0556_),
    .B(_0560_),
    .ZN(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1130_ (.A1(\writable[14] ),
    .A2(_0557_),
    .B(_0558_),
    .ZN(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1131_ (.A1(_0514_),
    .A2(_0556_),
    .B(_0561_),
    .ZN(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _1132_ (.A1(\writable[15] ),
    .A2(_0557_),
    .B(_0558_),
    .ZN(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _1133_ (.A1(_0516_),
    .A2(_0556_),
    .B(_0562_),
    .ZN(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1134_ (.D(_0000_),
    .CLK(clknet_2_1__leaf_wb_clk_i),
    .Q(\full_addr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1135_ (.D(_0001_),
    .CLK(clknet_2_1__leaf_wb_clk_i),
    .Q(\full_addr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1136_ (.D(_0002_),
    .CLK(clknet_2_1__leaf_wb_clk_i),
    .Q(\full_addr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1137_ (.D(_0003_),
    .CLK(clknet_2_1__leaf_wb_clk_i),
    .Q(\full_addr[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1138_ (.D(_0004_),
    .CLK(clknet_2_2__leaf_wb_clk_i),
    .Q(\full_addr[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _1139_ (.D(_0005_),
    .CLK(clknet_2_2__leaf_wb_clk_i),
    .Q(\full_addr[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1140_ (.D(_0006_),
    .CLK(clknet_2_2__leaf_wb_clk_i),
    .Q(\full_addr[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1141_ (.D(_0007_),
    .CLK(clknet_2_2__leaf_wb_clk_i),
    .Q(\full_addr[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1142_ (.D(_0008_),
    .CLK(clknet_2_0__leaf_wb_clk_i),
    .Q(\writable[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1143_ (.D(_0009_),
    .CLK(clknet_2_0__leaf_wb_clk_i),
    .Q(\writable[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1144_ (.D(_0010_),
    .CLK(clknet_2_0__leaf_wb_clk_i),
    .Q(\writable[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1145_ (.D(_0011_),
    .CLK(clknet_2_0__leaf_wb_clk_i),
    .Q(\writable[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1146_ (.D(_0012_),
    .CLK(clknet_2_3__leaf_wb_clk_i),
    .Q(\writable[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1147_ (.D(_0013_),
    .CLK(clknet_2_2__leaf_wb_clk_i),
    .Q(\writable[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1148_ (.D(_0014_),
    .CLK(clknet_2_2__leaf_wb_clk_i),
    .Q(\writable[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1149_ (.D(_0015_),
    .CLK(clknet_2_2__leaf_wb_clk_i),
    .Q(\writable[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1150_ (.D(_0016_),
    .CLK(clknet_2_3__leaf_wb_clk_i),
    .Q(\full_addr[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1151_ (.D(_0017_),
    .CLK(clknet_2_0__leaf_wb_clk_i),
    .Q(\full_addr[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1152_ (.D(_0018_),
    .CLK(clknet_2_3__leaf_wb_clk_i),
    .Q(\full_addr[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1153_ (.D(_0019_),
    .CLK(clknet_2_3__leaf_wb_clk_i),
    .Q(\full_addr[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1154_ (.D(_0020_),
    .CLK(clknet_2_3__leaf_wb_clk_i),
    .Q(\full_addr[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1155_ (.D(_0021_),
    .CLK(clknet_2_3__leaf_wb_clk_i),
    .Q(\full_addr[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1156_ (.D(_0022_),
    .CLK(clknet_2_3__leaf_wb_clk_i),
    .Q(\full_addr[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1157_ (.D(_0023_),
    .CLK(clknet_2_3__leaf_wb_clk_i),
    .Q(\full_addr[15] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1158_ (.D(_0024_),
    .CLK(clknet_2_1__leaf_wb_clk_i),
    .Q(\writable[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1159_ (.D(_0025_),
    .CLK(clknet_2_1__leaf_wb_clk_i),
    .Q(\writable[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1160_ (.D(_0026_),
    .CLK(clknet_2_1__leaf_wb_clk_i),
    .Q(\writable[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1161_ (.D(_0027_),
    .CLK(clknet_2_0__leaf_wb_clk_i),
    .Q(\writable[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1162_ (.D(_0028_),
    .CLK(clknet_2_3__leaf_wb_clk_i),
    .Q(\writable[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1163_ (.D(_0029_),
    .CLK(clknet_2_3__leaf_wb_clk_i),
    .Q(\writable[13] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1164_ (.D(_0030_),
    .CLK(clknet_2_2__leaf_wb_clk_i),
    .Q(\writable[14] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _1165_ (.D(_0031_),
    .CLK(clknet_2_3__leaf_wb_clk_i),
    .Q(\writable[15] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_wb_clk_i (.I(wb_clk_i),
    .Z(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_0__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_2_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_1__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_2_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_2__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_2_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_2_3__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_2_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input1 (.I(WEb_raw),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input10 (.I(cs_port[0]),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input11 (.I(cs_port[1]),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input12 (.I(cs_port[2]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input13 (.I(le_hi_act),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input14 (.I(le_lo_act),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input15 (.I(ram_end[0]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input16 (.I(ram_end[10]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input17 (.I(ram_end[11]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input18 (.I(ram_end[12]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input19 (.I(ram_end[13]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input2 (.I(bus_in[0]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input20 (.I(ram_end[14]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input21 (.I(ram_end[15]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input22 (.I(ram_end[1]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input23 (.I(ram_end[2]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input24 (.I(ram_end[3]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input25 (.I(ram_end[4]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input26 (.I(ram_end[5]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input27 (.I(ram_end[6]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input28 (.I(ram_end[7]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input29 (.I(ram_end[8]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(bus_in[1]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input30 (.I(ram_end[9]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input31 (.I(ram_start[0]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input32 (.I(ram_start[10]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input33 (.I(ram_start[11]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input34 (.I(ram_start[12]),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input35 (.I(ram_start[13]),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input36 (.I(ram_start[14]),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input37 (.I(ram_start[15]),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input38 (.I(ram_start[1]),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input39 (.I(ram_start[2]),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input4 (.I(bus_in[2]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input40 (.I(ram_start[3]),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input41 (.I(ram_start[4]),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input42 (.I(ram_start[5]),
    .Z(net42));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input43 (.I(ram_start[6]),
    .Z(net43));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input44 (.I(ram_start[7]),
    .Z(net44));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input45 (.I(ram_start[8]),
    .Z(net45));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input46 (.I(ram_start[9]),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input47 (.I(rom_enabled),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input48 (.I(rst),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(bus_in[3]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input6 (.I(bus_in[4]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input7 (.I(bus_in[5]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(bus_in[6]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input9 (.I(bus_in[7]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output49 (.I(net49),
    .Z(bus_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output50 (.I(net50),
    .Z(bus_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output51 (.I(net51),
    .Z(bus_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output52 (.I(net52),
    .Z(bus_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output53 (.I(net53),
    .Z(bus_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output54 (.I(net54),
    .Z(bus_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output55 (.I(net55),
    .Z(bus_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output56 (.I(net56),
    .Z(bus_out[7]));
endmodule

