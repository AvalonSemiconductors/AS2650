* NGSPICE file created from wrapped_as2650.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_1 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_2 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai33_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai33_1 A1 A2 A3 B1 B2 B3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyd_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyd_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_4 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_4 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

.subckt wrapped_as2650 io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ vdd vss wb_clk_i wb_rst_i
XFILLER_79_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6209__A2 _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7406__A1 _2656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7963_ _2537_ _3199_ _3200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6914_ _2212_ _2213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6425__I _1751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7894_ _2470_ _3131_ _3133_ _3134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_70_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7709__A2 _2939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6845_ _0804_ _0815_ _1832_ _2161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_126_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8382__A2 _3582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6776_ _2071_ _2094_ _2095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5196__A2 _4295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7590__B1 _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8515_ _1657_ _3484_ _3707_ _3711_ _3712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_104_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5727_ _1149_ _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4943__A2 _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8134__A2 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8446_ _3640_ _3641_ _3644_ _3645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5658_ as2650.pc\[8\] _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_108_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7893__A1 _2781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4609_ _4154_ _4190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8377_ _1407_ _3572_ _3577_ _2622_ _3578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_105_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5589_ _0589_ _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7328_ _1449_ _2586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_46_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4829__B _4408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7645__A1 _4307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7259_ _1280_ _2521_ _2522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_77_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6999__A3 _2289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4474__A4 _4054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7948__A2 _3185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output37_I net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6335__I _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7176__A3 _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6384__A1 as2650.stack\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7166__I _2437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8125__A2 _3343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6136__A1 _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6954__B _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5662__A3 _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4870__A1 _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6245__I _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4960_ _4299_ _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4622__A1 _4202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4891_ as2650.r0\[3\] _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6630_ _0751_ _1951_ _1952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6561_ _0847_ _0850_ _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8300_ _4393_ _4359_ _3502_ _3503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_5512_ _0912_ _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6127__A1 _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6492_ _1814_ _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6127__B2 _4015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8231_ as2650.stack\[7\]\[9\] _3440_ _3441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7875__A1 _2298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5443_ _0880_ _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4689__A1 _4267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8162_ _1747_ _0973_ _1750_ _3389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_86_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5374_ _0385_ _0807_ _0812_ _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_7113_ _2347_ _2384_ _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7627__A1 _2832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7627__B2 _2842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8093_ _2594_ _3324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7044_ _2322_ _2324_ _2326_ _2327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_101_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5102__A2 _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6850__A2 _1766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4861__A1 _4326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8995_ _0156_ clknet_leaf_12_wb_clk_i as2650.addr_buff\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7946_ _1121_ _3155_ _3184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7877_ _3111_ _3116_ _3117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_58_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5994__I _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8355__A2 _3532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8370__I _4097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6828_ _0735_ _2056_ _1848_ _2144_ _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5169__A2 _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6759_ _2040_ _2044_ _2077_ _2078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4916__A2 _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9118__D _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8107__A2 _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6118__A1 _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6118__B2 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7866__A1 _2779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6669__A2 _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8429_ _2933_ _3627_ _3628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5341__A2 _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7618__A1 _2863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8291__A1 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7094__A2 _2094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4852__A1 as2650.holding_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8972__CLK clknet_leaf_35_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4604__A1 _4147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8346__A2 _4374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8280__I _3483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4907__A2 _4104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7857__A1 _3097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5332__A2 _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7609__A1 _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8282__A1 _3461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7085__A2 _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8282__B2 _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5090_ _4213_ _0531_ _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4983__I _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8455__I _2668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6832__A2 _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4916__C _4203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8585__A2 _3125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7800_ _2781_ _3011_ _2789_ _3043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8780_ _0892_ _0899_ _3951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_65_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5992_ _1349_ _1350_ _0792_ _1259_ _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_75_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7731_ _2970_ _2974_ _2975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_80_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4943_ _0382_ _0383_ _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_127_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8190__I _3408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7662_ _1688_ _2907_ _2908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4874_ as2650.idx_ctrl\[1\] _4058_ _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8123__C _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6613_ _0839_ _1935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5556__C1 as2650.stack\[5\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7593_ _0915_ _2835_ _2837_ _2838_ _2839_ _2840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_119_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5020__A1 _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6544_ _1801_ _1867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5571__A2 _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7848__A1 _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6475_ _4286_ _4110_ _1798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7534__I _2781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8214_ _2177_ _3410_ _3427_ _3428_ _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5426_ _4361_ _4096_ _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5323__A2 _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8845__CLK clknet_leaf_69_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8145_ _1487_ _3283_ _0875_ _3373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5357_ _4222_ _0454_ _0777_ _0512_ _0779_ _0455_ _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_82_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5054__I _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8076_ _1619_ _3245_ _3308_ _2730_ _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_134_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5288_ _0432_ _0717_ _0722_ _0727_ _4204_ _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_82_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5087__A1 _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4893__I _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7027_ _4093_ _2311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8025__A1 _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8025__B2 _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7784__B1 _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8978_ _0139_ clknet_leaf_77_wb_clk_i as2650.r123_2\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7929_ _1120_ _3141_ _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8328__A2 _2787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5229__I _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7839__A1 _2685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7444__I _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5314__A2 _4318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6511__A1 _4186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7067__A2 _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8016__A1 _4005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8567__A2 _3460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6578__A1 _1878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4979__I2 as2650.r123_2\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5002__A1 _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8868__CLK clknet_leaf_46_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4590_ _4170_ _4171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_122_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7354__I _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6260_ _1627_ _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5305__A2 _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6502__A1 _4250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5211_ _0571_ _0573_ _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6191_ _1567_ _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5142_ _0319_ _0300_ _0398_ _0424_ _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_111_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5073_ _0512_ _0513_ _0514_ _0455_ _0454_ _0426_ _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XANTENNA__8007__A1 _3223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8118__C _3282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8901_ _0062_ clknet_3_7_0_wb_clk_i as2650.r123_2\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_8832_ _2518_ _3992_ as2650.psu\[4\] _3996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6569__A1 _4382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6569__B2 _4375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7230__A2 _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6033__A3 _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5975_ _1359_ _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8763_ _3922_ _3924_ _3925_ _3934_ _3935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_80_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4926_ _0369_ _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7714_ as2650.stack\[7\]\[5\] _1296_ _1045_ as2650.stack\[6\]\[5\] _0913_ _2959_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8694_ _2267_ _3869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7645_ _4307_ _2883_ _2891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4857_ _0300_ _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8730__A2 _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7692__C _2603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7576_ _1423_ _2824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4788_ _4367_ _4368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6741__A1 _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4888__I _4382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6527_ _1837_ _1839_ _1841_ _1849_ _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_88_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6458_ as2650.stack\[1\]\[4\] _1769_ _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5409_ as2650.r0\[3\] _0560_ _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9023__CLK clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6389_ _1689_ _1731_ _1732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8246__A1 _2419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7049__A2 _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8128_ _2482_ _0709_ _3357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8095__I _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8059_ _3258_ _2651_ _3292_ _1474_ _3243_ _3293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_9_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8970__D _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7439__I _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6980__A1 _4119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5783__A2 _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8721__A2 _3893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4798__I _4198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7174__I _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8485__A1 _3666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7902__I _3140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5422__I _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7460__A2 _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7349__I _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5223__A1 _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6253__I _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5760_ as2650.stack\[6\]\[13\] _1162_ _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_62_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6971__A1 _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5774__A2 _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4711_ _4291_ _4292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5691_ as2650.stack\[3\]\[10\] _1111_ _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7430_ _2311_ _0290_ _2265_ _2680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_124_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8712__A2 _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4642_ _4222_ _4223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6723__A1 _2037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5526__A2 _4136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7361_ _2615_ _2616_ _2617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9046__CLK clknet_leaf_40_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4573_ as2650.ins_reg\[2\] as2650.ins_reg\[3\] _4154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_144_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9100_ _0261_ clknet_leaf_50_wb_clk_i as2650.stack\[4\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6312_ _1670_ _1671_ _1673_ _1661_ _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_143_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7279__A2 _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7292_ _1260_ _1263_ _2551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9031_ _0192_ clknet_3_3_0_wb_clk_i as2650.cycle\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6243_ _1612_ _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6174_ _4288_ _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_48_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8129__B _2898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5125_ _0565_ _0566_ _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5056_ _0384_ _0389_ _0496_ _0497_ _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_66_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7203__A2 _2470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8815_ _4286_ _3979_ _3982_ _2519_ _3983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5214__A1 _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8746_ as2650.carry _3916_ _2534_ _3919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6962__A1 _1846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5958_ _4142_ _1343_ _1243_ _1344_ _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_90_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4909_ _4039_ _0352_ _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8677_ _3852_ _0591_ _3856_ _3857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5889_ _4109_ _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8164__B1 _3390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8703__A2 _2324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7628_ _2780_ _2872_ _2791_ _2875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5517__A2 _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4576__I0 as2650.holding_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7559_ _2740_ _2741_ _2806_ _2807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8467__A1 _1650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8219__A1 as2650.stack\[7\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_10_wb_clk_i_I clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6953__A1 _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5756__A2 _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9069__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6705__A1 _2023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_14_wb_clk_i clknet_3_3_0_wb_clk_i clknet_leaf_14_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_32_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6181__A2 _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8458__A1 _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8458__B2 _3461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6957__B _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7130__A1 _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8906__CLK clknet_leaf_62_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6449__S _1778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5692__A1 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4495__A2 _4075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6930_ _2209_ _2227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5995__A2 _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7197__A1 _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6861_ _2165_ _2174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8600_ _3596_ _3792_ _2620_ _3793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5812_ _1137_ _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6792_ _2072_ _2090_ _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6944__A1 _2067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8531_ _4097_ _3726_ _3727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5743_ _1143_ _1151_ _1159_ _0029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8697__A1 _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8462_ net52 _3630_ _3660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5674_ _1086_ _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7413_ _2375_ _2420_ _2663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_11_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4625_ as2650.psl\[3\] _4206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8393_ net31 _3523_ _3191_ _3594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8449__A1 _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7344_ _1249_ _2596_ _2599_ _2600_ _2601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_85_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4556_ _4007_ _4136_ _4137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4722__A3 _4137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7275_ _4285_ _2534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7121__A1 _4364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4487_ _4066_ _4067_ _4068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9014_ _0175_ clknet_leaf_15_wb_clk_i net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6226_ _1596_ _1597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6157_ as2650.r123_2\[3\]\[4\] _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5062__I _4191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5108_ _4267_ _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8621__A1 _3180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6088_ _1473_ _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5435__A1 _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5039_ _0479_ _0480_ _0463_ _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5738__A2 _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6935__A1 _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5946__B _4396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8729_ _0488_ _0509_ _0639_ _2096_ _3901_ _3902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__4946__B1 _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8137__B1 _3364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8688__A1 _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8041__C _2590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7360__A1 _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8929__CLK clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5910__A2 _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput20 net20 io_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_122_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7112__A1 _1859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput31 net31 io_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput42 net42 io_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_122_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7663__A2 _2908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6068__I _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8612__A1 _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7415__A2 _2276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7179__A1 _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5729__A2 _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4937__B1 _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8679__A1 _3851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5147__I _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5390_ _0761_ _0768_ _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_126_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5901__A2 _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4986__I net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7103__A1 _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4919__C _4367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7060_ _1057_ _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7654__A2 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6011_ _4243_ _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5665__A1 _4015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8603__A1 _3790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7406__A2 _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8603__B2 _3602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4935__B _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8193__I _3411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7962_ _2599_ _3194_ _3198_ _3199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6090__A1 _4127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6913_ _0888_ _1096_ _2212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_70_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7893_ _2781_ _3113_ _3132_ _2335_ _3133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_78_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6917__A1 _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6844_ _0797_ _1907_ _1965_ _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6775_ _2072_ _2090_ _2093_ _2094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_91_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7590__B2 as2650.stack\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8514_ _2732_ _3710_ _3711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5726_ _1148_ _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8445_ _3610_ _3642_ _3611_ _3643_ _3644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_5657_ _1086_ _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4608_ _4188_ _4189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8376_ _3571_ _3576_ _3577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5588_ _1017_ _1020_ _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4539_ as2650.cycle\[3\] _4120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7327_ _1257_ _2574_ _2552_ _1481_ _2585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_137_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7645__A2 _2883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7258_ _1282_ _2489_ _2521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6209_ _1283_ _1565_ _1556_ _1231_ _1583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_77_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7189_ _1421_ _2277_ _2460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_131_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8317__B _3518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5520__I _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6081__A1 _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6620__A3 _1935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4631__A2 as2650.ins_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6908__A1 _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7176__A4 _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8833__A1 _3952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5647__A1 _4297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4890_ _0333_ _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_36_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7572__A1 as2650.stack\[4\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7572__B2 as2650.stack\[5\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6261__I _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6560_ _1881_ _1882_ _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5583__B1 _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5511_ _0909_ _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6491_ _4196_ _1813_ _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7324__A1 _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6127__A2 _4392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8230_ _3435_ _3440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5442_ _0879_ _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4689__A2 _4269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5373_ _4179_ _0809_ _0811_ _4171_ _4348_ _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_8161_ _3387_ _3388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7112_ _1859_ _2376_ _2379_ _2383_ _2384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_8092_ _3277_ _0553_ _3323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7627__A2 _2834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8824__A1 _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5638__A1 _4163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7043_ _4195_ _1368_ _2325_ _2326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_86_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7820__I as2650.addr_buff\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4861__A2 _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8052__A2 _2767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8994_ _0155_ clknet_leaf_11_wb_clk_i as2650.addr_buff\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7945_ _2947_ _3174_ _3182_ _2600_ _3183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_70_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7876_ _3083_ _3067_ _3116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_23_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6827_ _1807_ _2142_ _2143_ _2144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7563__A1 _2809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6171__I _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6758_ _0517_ _2076_ _2045_ _2077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_104_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5709_ _1104_ _1133_ _1134_ _0020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7315__A1 _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6118__A2 _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8600__B _2620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6689_ _2006_ _2009_ _2010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_104_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8428_ _2887_ _3600_ _3627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_121_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7216__B _2484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8359_ net30 _3460_ _3560_ _3561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5515__I _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7618__A2 _2810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8815__A1 _4286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8815__B2 _2519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4852__A2 _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6054__A1 _4007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7554__A1 _2793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7554__B2 _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7306__A1 _2326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7857__A2 _2860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7609__A2 _2576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8806__A1 _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6256__I _1603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5160__I _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6045__A1 _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7793__A1 _2897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5991_ _4007_ _1370_ _1377_ _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_91_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7730_ _2886_ _2889_ _2932_ _2973_ _2974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
X_4942_ _4335_ _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_45_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7661_ _1683_ _2858_ _2907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7545__A1 _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4873_ _4367_ _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6612_ _4376_ _0470_ _1934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5556__B1 _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5556__C2 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7592_ as2650.stack\[5\]\[3\] _1177_ _0914_ _2839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6543_ as2650.r123_2\[2\]\[0\] _1865_ _1866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8420__B _3619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5308__B1 _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6474_ _0937_ _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5859__A1 _4032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8213_ _1640_ _3416_ _3417_ _3428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5425_ _4111_ _0353_ _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4531__A1 _4110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8144_ _3273_ _1475_ _3370_ _3371_ _3294_ _3372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5356_ _4264_ _0781_ _0794_ _4280_ _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_59_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8646__I net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8273__A2 _2546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7076__A3 _2352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8075_ _3297_ _3306_ _3307_ _3308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5287_ _0726_ _4247_ _4252_ _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5087__A2 _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7026_ _4268_ _2302_ _2310_ _0161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8025__A2 _3258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5070__I _4275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6036__A1 _4080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8977_ _0138_ clknet_leaf_58_wb_clk_i as2650.stack\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7784__A1 _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7784__B2 _2312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4598__A1 _4178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7928_ _2640_ _3166_ _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7859_ _1256_ _3099_ _4293_ _3100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_93_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4770__A1 _4192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4522__A1 as2650.cycle\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7067__A3 _2314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_39_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_39_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6275__A1 _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8016__A2 _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6027__A1 _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7775__A1 _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4589__A1 _4027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4979__I3 as2650.r123_2\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5538__B1 _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5002__A2 _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5305__A3 _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6502__A2 _1824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5156__I3 as2650.r123_2\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5210_ _0614_ _0621_ _0650_ _4281_ _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_6190_ _4044_ _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5141_ _0530_ _0532_ _0534_ _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6266__A1 _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5072_ _0425_ _0444_ _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_69_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8900_ _0061_ clknet_leaf_74_wb_clk_i as2650.r123_2\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8831_ _2533_ _3995_ _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_92_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7766__A1 _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6569__A2 _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8762_ _3927_ _3929_ _3931_ _3933_ _3934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5974_ _1347_ _1357_ _1360_ _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7713_ as2650.stack\[4\]\[5\] _1192_ _2956_ as2650.stack\[5\]\[5\] _2958_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4925_ _0368_ _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7518__A1 _2761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8693_ _2431_ _1576_ _3868_ _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7644_ _2887_ _2889_ _2890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4856_ _4383_ _4385_ _4387_ _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XFILLER_20_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7575_ _2676_ _2823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4787_ _4024_ _4366_ _4367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6526_ _1842_ _1824_ _1844_ _1848_ _1849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__4752__A1 _4232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6457_ _1629_ _1774_ _1784_ _0118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8962__CLK clknet_leaf_77_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4504__A1 _4079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5408_ _0843_ _0844_ _0846_ _0763_ _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_88_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6388_ _1714_ _1731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8127_ _3338_ _3356_ _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_138_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5339_ _0599_ _0705_ _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6257__A1 _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6257__B2 as2650.stack\[5\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8058_ _2336_ _4400_ _3291_ _3292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_25_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4807__A2 _4386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7009_ as2650.addr_buff\[2\] _2298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7757__B2 as2650.stack\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6980__A2 _4118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4991__A1 _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8182__A1 _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4743__A1 _4138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8485__A2 _3680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7404__B _2590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8237__A2 _3440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7190__I _2460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6248__A1 _1615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8219__C _3408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5471__A2 _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7748__A1 _2546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5223__A2 _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6420__A1 _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6971__A2 _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4710_ _4037_ _4291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5690_ _1117_ _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8173__A1 _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4989__I _4226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4641_ _4221_ _4222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_129_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7920__A1 _2736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6723__A2 _2042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8985__CLK clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5526__A3 _4412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4734__A1 _4309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7360_ _1064_ _2257_ _2616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4572_ _4152_ _4153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_116_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6311_ as2650.stack\[4\]\[1\] _1672_ _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__8476__A2 _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7291_ _4079_ _2550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9030_ _0191_ clknet_leaf_15_wb_clk_i as2650.cycle\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_118_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6242_ as2650.pc\[1\] _1612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8228__A2 _3438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6173_ _4035_ _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_124_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6239__A1 _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5124_ _4381_ _0368_ _0466_ _4229_ _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7987__A1 _2530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5055_ _0395_ _0345_ _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7968__C _2685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7739__A1 _2576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8145__B _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8814_ _2504_ _3911_ _3974_ _3981_ _3982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_111_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5214__A2 _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8745_ _3917_ _3918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_111_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5957_ _4143_ _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6962__A2 _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4908_ _0350_ _0351_ _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8676_ _1635_ _3843_ _3856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5888_ _1282_ _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8164__A1 _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8164__B2 as2650.stack\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7627_ _2832_ _2834_ _2841_ _2842_ _2873_ _2874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4839_ _4418_ _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7911__A1 _3147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7275__I _4285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7558_ _4391_ _4233_ _2806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4576__I1 _4153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6112__C _1497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6509_ _1802_ _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7489_ _1613_ _2703_ _2738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_122_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8039__C _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7978__A1 _2464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8858__CLK clknet_leaf_58_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6953__A2 _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8155__A1 _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6705__A2 _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4716__A1 _4166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8458__A2 _3484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_54_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_99_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7130__A2 _2401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5141__A1 _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9052__D _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5692__A2 _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7969__A1 _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8091__B1 _3312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7433__A3 _2666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6264__I _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6860_ _1611_ _2167_ _2173_ _0132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7197__A2 _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5811_ _1207_ _1198_ _1208_ _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6791_ _2072_ _2090_ _2109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8530_ _1488_ _0780_ _3726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4955__A1 _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5742_ as2650.stack\[5\]\[14\] _1149_ _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8146__A1 _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8461_ _3625_ _3657_ _3658_ _3659_ _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5673_ _1102_ _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8697__A2 _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5608__I _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7412_ _1487_ _2535_ _2660_ _2662_ _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_50_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4624_ _4204_ _4205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8392_ _1729_ _3490_ _3592_ _2572_ _3593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_124_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7343_ _2466_ _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4555_ _4024_ _4107_ _4117_ _4135_ _4136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_85_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7274_ _2531_ _2378_ _2533_ _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_132_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4486_ _4041_ _4067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9013_ _0174_ clknet_leaf_14_wb_clk_i net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5132__A1 _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6225_ as2650.pc\[0\] _1596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7979__B _3214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6880__A1 _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5683__A2 _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6156_ _1537_ _0064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5107_ _4369_ _0548_ _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6087_ _1358_ _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_39_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5435__A2 _4299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5038_ _0463_ _0479_ _0480_ _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_38_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6174__I _4288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8385__A1 _2897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6935__A2 _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6989_ _4293_ _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8728_ _0407_ _0413_ _0628_ _0510_ _3900_ _3901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_55_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4946__B2 _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8137__A1 _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8137__B2 _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8659_ _3830_ _3836_ _3842_ _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4422__I _4002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6699__A1 _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7360__A2 _2257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput21 net21 io_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_122_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput32 net32 io_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput43 net43 io_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__5123__A1 _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6871__A1 _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8073__B1 _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5426__A2 _4096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6623__A1 _1941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9036__CLK clknet_leaf_40_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6084__I _4285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7179__A2 _2449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8128__A1 _2482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4937__B2 _4316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8679__A2 _3857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8300__A1 _4393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7103__A2 _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6259__I _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5163__I _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5665__A2 _4288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6862__A1 _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6010_ _1393_ _1396_ _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input3_I io_in[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8603__A2 _3793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7961_ _4095_ _2861_ _2708_ _1353_ _3198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_94_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6912_ as2650.r123_2\[0\]\[0\] _2208_ _2211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6090__A2 _1475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7892_ _2891_ _3125_ _3132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8367__A1 _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6843_ _0781_ _1810_ _2056_ _2158_ _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_63_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8423__B _3622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6917__A2 _2213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6774_ _2006_ _2009_ _2091_ _2092_ _2093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_51_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8119__A1 _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7590__A2 _2836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8513_ _1656_ _3491_ _3709_ _3654_ _3042_ _3710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5725_ _1145_ _1147_ _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8444_ _0539_ _0552_ _3643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5656_ _1085_ _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4607_ _4187_ _4188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8375_ _1484_ _0452_ _3575_ _3576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_5587_ _0916_ _1018_ _1019_ _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_117_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7326_ _1230_ _1237_ _2584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4538_ as2650.cycle\[1\] _4119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_105_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6169__I _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7257_ _2520_ _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4469_ as2650.cycle\[5\] _4050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6208_ _1231_ _1555_ _1549_ _1581_ _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_104_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6853__A1 _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7188_ _2458_ _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__9059__CLK clknet_leaf_40_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6139_ _1522_ _1524_ _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_86_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7802__B1 _3019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8358__A1 _3461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4919__A1 _4258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5592__A1 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8530__A1 _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6136__A3 _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5895__A2 _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7097__A1 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8833__A2 _3991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6844__A1 _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5647__A2 _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8349__A1 _3549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7638__I _2883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7021__A1 _2307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5510_ _0881_ _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6490_ _1812_ _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7324__A2 _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5441_ _0875_ _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5335__B2 _4316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7373__I _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8160_ _1602_ _1160_ _3387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5372_ _0641_ _0716_ _0810_ _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7111_ _2258_ _2382_ _2383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7088__A1 _4412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8091_ _1628_ _3276_ _3312_ _3322_ _2639_ _0214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__8824__A2 _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5638__A2 _4089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7042_ _2283_ _2325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8588__A1 _3772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8588__B2 _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8993_ _0154_ clknet_leaf_69_wb_clk_i as2650.r123_2\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8919__CLK clknet_leaf_33_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7944_ _2796_ _3168_ _3181_ _1256_ _1354_ _3182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_23_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5810__A2 _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7875_ _2298_ _3114_ _3115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_36_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7548__I _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6826_ _0709_ _1918_ _2143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7563__A2 _2810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8760__A1 _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7992__B _4260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6757_ _1936_ _2076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5708_ as2650.stack\[3\]\[12\] _1111_ _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_137_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6688_ _1927_ _2007_ _2008_ _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__8512__A1 _3326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7315__A2 _2539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8427_ _2580_ _3626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5326__A1 as2650.r0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5639_ _4080_ _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7283__I _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4700__I _4135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8358_ _3461_ _3557_ _3559_ _3485_ _3560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_2_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7079__A1 _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7309_ _2481_ _2344_ _2566_ _2567_ _2568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_8289_ _1248_ _1547_ _3492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_137_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6826__A1 _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7232__B _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5531__I _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6054__A2 _1440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5801__A2 _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7458__I _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6362__I _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7554__A2 _2795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8503__A1 net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7306__A2 _2564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5317__A1 _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7193__I _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8267__B1 _3470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7609__A3 _2855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8806__A2 _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7490__A1 _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5441__I _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6045__A2 _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5990_ _0521_ _1374_ _1376_ _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_91_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4941_ _0382_ _0383_ _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_79_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5089__S _4012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7660_ _2898_ _2903_ _2904_ _2905_ _2906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_127_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4872_ _0315_ _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7545__A2 _2736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8742__A1 _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6611_ _1883_ _1899_ _1932_ _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7591_ as2650.stack\[7\]\[3\] _2697_ _1047_ as2650.stack\[6\]\[3\] _2836_ as2650.stack\[4\]\[3\]
+ _2838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
X_6542_ _1864_ _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_9_wb_clk_i clknet_3_2_0_wb_clk_i clknet_leaf_9_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7317__B _2574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5308__A1 _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5308__B2 _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6473_ _1654_ _1774_ _1796_ _0122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5616__I _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5859__A2 _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8212_ as2650.stack\[7\]\[4\] _3413_ _3427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5424_ _4111_ _4086_ _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8143_ _3340_ _0797_ _3324_ _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5355_ _4200_ _0791_ _0793_ _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4531__A2 _4111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6808__A1 _1962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8074_ _1568_ _0357_ _3263_ _2014_ _3243_ _3307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_101_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5286_ _0725_ _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_87_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8148__B _3375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7025_ _1584_ _2304_ _2310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6447__I _4377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7481__A1 _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6036__A2 _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8976_ _0137_ clknet_leaf_58_wb_clk_i as2650.stack\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5244__B1 _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7784__A2 _2804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8891__CLK clknet_leaf_51_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4598__A2 _4170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7927_ _1122_ _2686_ _3165_ _3166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_58_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6182__I _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7858_ _2743_ _3098_ _3099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6809_ _2121_ _2118_ _2126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7789_ _1372_ _0595_ _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_71_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4770__A2 _4239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4430__I _4010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7472__A1 _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5261__I _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7224__A1 _2488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6027__A2 _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8421__B1 _3620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8505__C _3626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4589__A2 _4070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7188__I _2458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9055__D _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5140_ _0535_ _0580_ _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_123_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5071_ _0491_ _0448_ _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5104__C _4204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8830_ _3992_ _3993_ _3994_ _3995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8415__C _2626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5777__A1 _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8761_ _1265_ _1464_ _2480_ _3932_ _3933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_5973_ _1359_ _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7712_ as2650.stack\[0\]\[5\] _1192_ _2956_ as2650.stack\[1\]\[5\] _0921_ _2957_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_4924_ _0367_ _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8692_ _2303_ _1573_ _3868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8715__A1 as2650.psl\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7643_ _2844_ _2848_ _2888_ _2889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_61_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5529__A1 _4308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4855_ _4165_ _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7574_ _0914_ _2816_ _2817_ _2821_ _2822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_4786_ _4362_ _4364_ _4365_ _4366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_119_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6525_ _1847_ _1095_ _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5346__I _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6456_ as2650.stack\[1\]\[3\] _1768_ _1783_ _1773_ _1784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_118_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5407_ _0564_ _0525_ _0845_ _0665_ _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5701__A1 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4504__A2 _4084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7561__I _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6387_ _1727_ _1722_ _1728_ _1730_ _0102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8126_ _3355_ _1734_ _3244_ _3356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5338_ _0715_ _0776_ _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_130_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8057_ _1401_ _1396_ _3290_ _2603_ _3291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5269_ _0708_ _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7008_ _2297_ _0156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7510__B _2758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8959_ _0120_ clknet_leaf_47_wb_clk_i as2650.stack\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4425__I _4005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6193__A1 _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8060__C _2639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4743__A2 _4283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6087__I _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7996__A2 _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7748__A2 _2991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5759__A1 _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5223__A3 _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7646__I _2891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4640_ _4211_ _4216_ _4220_ _4221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__6184__A1 _4032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7920__A2 _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4571_ _4148_ _4149_ _4150_ _4151_ _4018_ _4019_ _4152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__4734__A2 _4314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5931__A1 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6310_ _1664_ _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7290_ _2341_ _2548_ _2549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6241_ _1610_ _1611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7684__A1 _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4498__A1 _4072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6172_ _1548_ _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5123_ _0563_ _0564_ _0368_ _0465_ _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_58_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5054_ _0407_ _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_22_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9092__CLK clknet_leaf_26_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8813_ _1264_ _3975_ _3980_ _3981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_0_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5956_ _1342_ _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_8744_ _3913_ _3914_ _3916_ _3917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4907_ _4063_ _4104_ _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8675_ _3851_ _3854_ _3855_ _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_142_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7556__I _2803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5887_ _1281_ _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7626_ _2856_ _2871_ _2872_ _2873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4838_ _4376_ _4188_ _4321_ _4417_ _4418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_14_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7557_ net7 _4384_ _2805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_105_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5076__I _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4769_ _4326_ _4191_ _4349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6508_ _4272_ _1810_ _1830_ _1807_ _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_119_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7488_ _2735_ _2736_ _2737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6439_ as2650.stack\[1\]\[0\] _1769_ _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7291__I _4079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7427__A1 _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8109_ _3324_ _2096_ _3339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9089_ _0250_ clknet_leaf_26_wb_clk_i net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5989__A1 _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_4_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8055__C _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8071__B _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4964__A2 _4191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8155__A2 _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8297__I _2559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7666__A1 _2910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7418__A1 _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_23_wb_clk_i clknet_opt_3_1_wb_clk_i clknet_leaf_23_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_132_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7969__A2 _2731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8091__A1 _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7197__A3 _2456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5810_ as2650.stack\[1\]\[12\] _1201_ _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_63_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8952__CLK clknet_leaf_59_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6790_ as2650.r123_2\[2\]\[5\] _2069_ _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5601__B1 _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5741_ _1138_ _1151_ _1158_ _0028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4955__A2 _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6280__I _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8460_ _1294_ _3659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5672_ _1088_ _1090_ _1098_ as2650.r123_2\[0\]\[0\] _1101_ _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_124_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8697__A3 _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7411_ _1039_ _2374_ _2661_ net4 _0861_ _2662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_15_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4623_ _4203_ _4204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8391_ _3581_ _3584_ _3591_ _3592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4707__A2 _4284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7342_ _2598_ _2599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4554_ _4134_ _4135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5380__A2 _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7657__A1 _2900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7273_ _2532_ _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4485_ _4065_ _4066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_9012_ _0173_ clknet_leaf_4_wb_clk_i as2650.r123\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6224_ _1594_ _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7409__A1 _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8606__B1 _3798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6155_ as2650.r123_2\[3\]\[3\] _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7979__C _2335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5106_ _0518_ _4378_ _0547_ _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8082__A1 _4206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6086_ _1470_ _1472_ _0059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5037_ _0474_ _0475_ _0477_ _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_73_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5435__A3 _4300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4643__A1 _4207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8670__I _3835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8385__A2 _3564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6988_ _2262_ _2264_ _2266_ _2278_ _2279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__8603__C _2458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8727_ _3891_ _3894_ _3899_ _3900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7286__I _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5939_ _0625_ _0629_ _1325_ _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8137__A2 _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6190__I _4044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4703__I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6148__A1 _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7219__C _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8658_ _3838_ _3262_ _3839_ _3841_ _3842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_90_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7896__A1 _2779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7609_ _1336_ _2576_ _2855_ _2856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6699__A2 _1973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8589_ _1114_ _3490_ _3782_ _3461_ _3783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_31_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5371__A2 _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput11 net11 io_oeb[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_134_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput22 net22 io_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_134_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput33 net52 io_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput44 net44 io_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_107_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4882__A1 _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4882__B2 _4356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8073__A1 _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8073__B2 _3305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8066__B _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8975__CLK clknet_leaf_59_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8376__A2 _3576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6387__A1 _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8513__C _3042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4937__A2 _4413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8128__A2 _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4613__I _4075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7887__A1 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5362__A2 _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7639__A1 _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5444__I _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8300__A2 _4359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7103__A3 _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5114__A2 _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6311__A1 as2650.stack\[4\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8064__A1 _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7960_ _1135_ _3196_ _3197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6911_ _2209_ _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7891_ _3039_ _3115_ _3117_ _3029_ _2600_ _3130_ _3131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__8367__A2 _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6842_ _1844_ _2157_ _2158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6378__A1 _1615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8423__C _3485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6773_ _2028_ _2029_ _2053_ _2092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8119__A2 _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8512_ _3326_ _3700_ _3708_ _3709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5724_ _1146_ _0988_ _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7327__B1 _2552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7878__A1 as2650.pc\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8443_ _0538_ _0552_ _3642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5655_ _1044_ _1048_ _1084_ _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_108_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4606_ _4148_ _4187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8374_ _3549_ _3573_ _3574_ _3575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8848__CLK clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5586_ as2650.stack\[7\]\[13\] _0977_ _0900_ as2650.stack\[6\]\[13\] _1019_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_117_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7325_ _2344_ _2567_ _2582_ _2583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_116_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4537_ _4033_ _4118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_11_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5105__A2 _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7256_ _0490_ _2519_ _2501_ _2520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_104_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4468_ _4043_ _4049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_131_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6207_ _1580_ _1544_ _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_63_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8998__CLK clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6853__A2 _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7187_ _2427_ _2410_ _2458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8055__A1 _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6138_ _1518_ _1523_ _1266_ _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6185__I _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7802__A1 _2832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7802__B2 _2842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6069_ _0405_ _1250_ _1449_ _1455_ _1345_ _4196_ _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai33_1
XTAP_3227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4616__A1 _4082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4634__S _4013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6369__A1 as2650.stack\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7566__B1 _2812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4919__A2 _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5041__A1 _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4433__I _4013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8530__A2 _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7097__A2 _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9003__CLK clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5647__A3 _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6095__I _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4608__I _4188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7021__A2 _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5583__A2 _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6780__A1 _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7324__A3 _2560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5440_ _0877_ _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5335__A2 _4413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5371_ _0799_ _0641_ _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5174__I _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7110_ _2380_ _2381_ _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7088__A2 _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8090_ _2303_ _3264_ _3259_ _3319_ _3321_ _3322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_99_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8824__A3 _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7041_ _1442_ _2323_ _2324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5638__A3 _4074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5902__I _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8037__A1 _3271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6599__A1 _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8992_ _0153_ clknet_leaf_46_wb_clk_i as2650.r123_2\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_94_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout54_I net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7943_ _2905_ _3180_ _3181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7829__I _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7874_ _3062_ _3097_ _3065_ _3114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_63_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_7_0_wb_clk_i clknet_0_wb_clk_i clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_6825_ _1810_ _2141_ _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8760__A2 _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7992__C _2656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6756_ _2073_ _2074_ _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5707_ _1132_ _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6687_ _1930_ _1959_ _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_52_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8426_ _3488_ _3625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5638_ _4163_ _4089_ _4074_ _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_30_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9026__CLK clknet_leaf_17_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8357_ _1623_ _3558_ _3559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5569_ as2650.stack\[0\]\[12\] _0953_ _0972_ as2650.stack\[1\]\[12\] _1003_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_88_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7308_ _1578_ _1433_ _2567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7079__A2 _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8288_ _3479_ _3491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8609__B _3485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6826__A2 _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7239_ _2505_ _2506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_63_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_69_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7232__C _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6129__B _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6054__A3 _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output35_I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8063__C _2547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8200__A1 _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5014__A1 _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5014__B2 _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5565__A2 _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7474__I _2430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5317__A2 _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8267__A1 _3464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8267__B2 _2256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4828__A1 _4377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8019__A1 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7242__A2 _2507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5253__A1 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4940_ as2650.holding_reg\[3\] _0345_ _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_45_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4871_ _0298_ _0314_ _4146_ _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5005__A1 _4265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8742__A2 _2550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6610_ _1885_ _1898_ _1932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7590_ as2650.stack\[0\]\[3\] _2836_ _2695_ as2650.stack\[1\]\[3\] _2837_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__5556__A2 _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6541_ _1801_ _1863_ _1864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__9049__CLK clknet_leaf_40_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4801__I as2650.r0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5308__A2 _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6472_ as2650.stack\[1\]\[7\] _1768_ _1795_ _1773_ _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__6505__A1 _4224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5423_ _4110_ _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8211_ _1727_ _3419_ _3426_ _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_127_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8258__A1 _2620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8142_ _2623_ _0781_ _3370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5354_ _0792_ _4200_ _4258_ _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6808__A2 _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8073_ _2299_ _3264_ _3259_ _3305_ _3306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5285_ _0724_ _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_138_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7024_ _4266_ _2302_ _2309_ _0160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7481__A2 _2686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8975_ _0136_ clknet_leaf_59_wb_clk_i as2650.stack\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5244__B2 _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7926_ _2894_ _3142_ _3163_ _3164_ _2684_ _3165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_93_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6992__A1 _4035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7857_ _3097_ _2860_ _3098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5079__I _4019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8733__A2 _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6808_ _1962_ _2107_ _2108_ _2125_ _0128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4912__S _4238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5547__A2 _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6744__A1 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7788_ _1794_ _3030_ _3031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6739_ _1409_ _1910_ _2057_ _1836_ _2058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_20_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4711__I _4291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6131__C _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8409_ _1411_ _3603_ _3507_ _3608_ _3609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__8249__A1 _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8339__B _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7472__A2 _2713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5483__A1 _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8421__A1 _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7224__A2 _2491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8421__B2 _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7775__A3 _3017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6983__A1 _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5786__A2 _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8802__B _3969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_48_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__8724__A2 _4353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5538__A2 _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8488__A1 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7160__A1 _4070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4777__B _4276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7463__A2 _2712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5070_ _4275_ _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_78_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5474__A1 _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6283__I _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8760_ _1500_ _1259_ _2883_ _3932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5972_ _1358_ _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5777__A2 _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7711_ _1175_ _2956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4923_ as2650.r123\[0\]\[2\] as2650.r123_2\[0\]\[2\] _4008_ _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8691_ _3851_ _3866_ _3867_ _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_90_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8715__A2 _3882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7642_ _2845_ _2888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4854_ _0297_ _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4785_ as2650.idx_ctrl\[1\] as2650.idx_ctrl\[0\] _4365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7573_ _0922_ _2818_ _2820_ _2821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__5627__I _4118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6524_ _0641_ _4127_ _4132_ _1846_ _1847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_105_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4752__A3 _4236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7151__A1 _2343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6455_ _1684_ _1782_ _1783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5406_ _0765_ _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6386_ _1729_ _1718_ _1719_ _1730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5701__A2 _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8125_ _3339_ _3343_ _3353_ _3354_ _3355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5337_ _0680_ _0703_ _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8651__A1 _3223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5268_ _0443_ _0600_ _0704_ _0550_ _0707_ _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__7454__A2 _2265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8056_ _3281_ _0355_ _3289_ _1395_ _3290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_9_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5465__A1 _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7007_ _2296_ _1572_ _2294_ _2297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_87_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5199_ _4193_ _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__8606__C _2437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7206__A2 _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7289__I _4081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4706__I as2650.halted vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8958_ _0119_ clknet_leaf_47_wb_clk_i as2650.stack\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7909_ as2650.pc\[10\] _1491_ _3148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8889_ _0050_ clknet_leaf_64_wb_clk_i as2650.stack\[1\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6717__A1 _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7914__B1 _3151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4991__A3 _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7390__A1 _4364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6193__A2 _1563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5537__I _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4441__I _4021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7142__A1 _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7752__I _2760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8069__B _3301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5272__I _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7701__B _2869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7996__A3 _3225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7199__I _2469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5208__A1 _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5759__A2 _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6956__A1 _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4806__I1 as2650.r123\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7148__B _2419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4570_ as2650.r123\[2\]\[0\] as2650.r123_2\[2\]\[0\] _4009_ _4151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7133__A1 _2286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6240_ _4230_ _1610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8881__CLK clknet_leaf_47_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4498__A2 _4078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6171_ _1547_ _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5122_ as2650.r0\[1\] _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5447__A1 _4311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5053_ _0494_ _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4670__A2 _4250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8812_ _2374_ _3976_ _3980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8743_ _3880_ _3915_ _3916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5955_ _1341_ _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4906_ _4143_ _4099_ _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8674_ net44 _3846_ _3855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5886_ _0604_ _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_16_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7058__B _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7625_ _2647_ _2834_ _2849_ _2472_ _2537_ _2872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_4837_ _4416_ _4417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7556_ _2803_ _2804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5922__A2 _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6897__B _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4768_ _4140_ _4168_ _4348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6507_ _1588_ _1816_ _1828_ _1829_ _1830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_119_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7487_ _2538_ _2736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4699_ _4273_ _4280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6438_ _1767_ _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6369_ as2650.stack\[3\]\[0\] _1715_ _1716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8624__A1 _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7427__A2 _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8108_ _2532_ _3338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9088_ _0249_ clknet_leaf_26_wb_clk_i net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8624__B2 _2485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5438__A1 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8039_ _3271_ _4279_ _3272_ _3273_ _3274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_29_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5989__A2 _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6938__A1 _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5610__A1 _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6166__A2 _4054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7363__A1 _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8560__B1 _3754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5913__A2 _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6098__I _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8615__A1 net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7418__A2 _4081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8091__A2 _3276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7197__A4 _2467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5601__A1 as2650.stack\[3\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5740_ as2650.stack\[5\]\[13\] _1149_ _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5671_ _0933_ _1099_ _1100_ _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8697__A4 _2314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7410_ _2374_ _2658_ _2661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4622_ _4202_ _4197_ _4203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8390_ _1631_ _2586_ _3585_ _3590_ _3591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_102_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7606__B _2606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7341_ _1577_ _2353_ _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4553_ _4017_ _4133_ _4134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7106__A1 _4307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4484_ _4064_ _4065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7272_ _1293_ _2532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9011_ _0172_ clknet_leaf_0_wb_clk_i as2650.r123\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6223_ _1593_ _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8606__A1 _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6154_ _1536_ _0063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7409__A2 _2657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8606__B2 _2668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8437__B _4060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5105_ _4240_ _0346_ _0546_ _4198_ _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8082__A2 _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6085_ _1375_ _1468_ _1471_ _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5036_ _0478_ _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5435__A4 _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4643__A2 _4223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5840__A1 _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6987_ _2267_ _1062_ _2274_ _2277_ _2278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_53_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7593__A1 _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8726_ _0315_ _3893_ _3897_ _3898_ _3899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_107_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5938_ _0647_ _0639_ _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8657_ _1589_ _3840_ _3841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7345__A1 _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6148__A2 _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5869_ _1258_ _1260_ _1263_ _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7608_ _2850_ _2853_ _2854_ _2855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_8588_ _3772_ _3776_ _3781_ _1360_ _3782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_124_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7539_ _2785_ _2786_ _2787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_119_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput12 net12 io_oeb[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput23 net23 io_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_135_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput34 net34 io_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput45 net45 io_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_122_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4882__A2 _4389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8073__A2 _3264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5831__A1 _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7477__I _2683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7887__A2 _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9082__CLK clknet_leaf_25_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7639__A2 _2884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8064__A2 _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6075__A1 _4260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6910_ _0939_ _1096_ _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7890_ _2843_ _3125_ _3112_ _2796_ _3129_ _3130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_35_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8367__A3 _3567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6841_ _1039_ _1908_ _2156_ _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_78_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7387__I _2639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6291__I as2650.pc\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5586__B1 _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6772_ _2028_ _2053_ _2091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8511_ _2558_ _2862_ _3708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5723_ _1043_ _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7327__A1 _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7327__B2 _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8442_ _3639_ _0586_ _3641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7878__A2 _2987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5654_ _1083_ _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4605_ _4147_ _4159_ _4185_ _4186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_8373_ _0348_ _0330_ _3574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6550__A2 _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5585_ as2650.stack\[4\]\[13\] _0971_ _0918_ as2650.stack\[5\]\[13\] _1018_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8011__I _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7324_ _2428_ _2440_ _2560_ _2581_ _2582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_105_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4536_ _4109_ _4112_ _4116_ _4117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_144_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7255_ _1635_ _2517_ _2518_ _2519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_4467_ _4047_ _4048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_131_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6206_ _1442_ _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7186_ _1064_ _2456_ _2457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6853__A3 _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_59_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6137_ _1499_ _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8055__A2 _3262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6066__A1 _4310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7802__A2 _3011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6068_ _1454_ _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_39_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4616__A2 _4112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5019_ _4302_ _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6081__A4 _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7566__A1 _2735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7566__B2 _2813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4714__I _4115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5041__A2 _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8709_ _1266_ _1280_ _3883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7869__A2 _2686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5545__I _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4552__A1 _4125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8818__A1 _2515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8818__B2 _4206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8942__CLK clknet_leaf_43_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8046__A2 _4355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7557__A1 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4624__I _4204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7309__A1 _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4543__A1 _4118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8809__A1 _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5370_ _0802_ _0808_ _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_141_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6296__A1 _1654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7040_ _4035_ _1562_ _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6286__I _1650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8037__A2 _4272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6048__A1 _4007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8991_ _0152_ clknet_leaf_68_wb_clk_i as2650.r123_2\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8715__B _3888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7942_ as2650.addr_buff\[4\] _2803_ _3180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7873_ _3112_ _3113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_51_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6824_ _0712_ _1971_ _2140_ _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6220__A1 _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6755_ _1987_ _2048_ _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8450__B _3579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5706_ _1130_ _1090_ _1098_ as2650.r123_2\[0\]\[4\] _1131_ _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_91_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6686_ _1930_ _1959_ _2007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_17_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8425_ _3595_ _3624_ _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5637_ _1052_ _1066_ _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6523__A2 _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7720__A1 _2591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8965__CLK clknet_leaf_76_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7720__B2 _2931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8356_ _1359_ _2490_ _2485_ _3558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_128_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5568_ as2650.stack\[2\]\[12\] _0920_ _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7307_ _4056_ _2540_ _2560_ _2565_ _2566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_137_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4519_ _4062_ _4099_ _4100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8287_ _3483_ _3490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5499_ _4108_ _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6287__A1 _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7238_ _1401_ _1355_ _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_137_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6196__I _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4709__I _4289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7169_ _2341_ _1552_ _2439_ net54 _2440_ _2441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_115_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6039__A1 _4260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5262__A2 _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6145__B _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output28_I net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5014__A2 _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8998__D _0159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4773__A1 _4331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7011__I0 _2298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4525__A1 _4039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7475__B1 _2722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9120__CLK clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7490__A3 _2738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7778__A1 _1650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5253__A2 _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4870_ _0299_ _0295_ _0311_ _0313_ _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5005__A2 _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8742__A3 _2677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6753__A2 _2052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8988__CLK clknet_leaf_69_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7950__A1 _2760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6540_ _1520_ _1862_ _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6471_ _1794_ _1782_ _1795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8210_ as2650.stack\[7\]\[3\] _3424_ _3425_ _3409_ _3426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__4516__A1 _4093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5422_ _0528_ _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8141_ _3338_ _3369_ _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8258__A2 _2713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5353_ _4210_ _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8072_ _1385_ _1495_ _3302_ _3304_ _3305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_87_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5284_ _0723_ _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_82_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7023_ _1283_ _2304_ _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8974_ _0135_ clknet_leaf_57_wb_clk_i as2650.stack\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6441__A1 _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7925_ _0994_ _2690_ _3157_ _2689_ _2687_ _3164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_58_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6992__A2 _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7856_ as2650.addr_buff\[1\] _3097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_24_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6807_ _2071_ _2124_ _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7787_ _1737_ _2984_ _3030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__7575__I _2676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7941__A1 _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4999_ _0415_ _4200_ _4370_ _0441_ _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6744__A2 _1966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4755__A1 _4178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6738_ _0543_ _1823_ _2057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6669_ _0417_ _0845_ _1990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5095__I _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8408_ _3603_ _3607_ _3608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8249__A2 _2666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8339_ _0321_ _0326_ _0347_ _3541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5180__A1 _4135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4867__C _4348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6680__A1 _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8421__A2 _3525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8074__C _3243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5235__A2 _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6432__A1 _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6983__A2 _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8185__A1 _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7485__I _2733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7932__A1 _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6735__A2 _2054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4902__I _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_17_wb_clk_i clknet_opt_1_0_wb_clk_i clknet_leaf_17_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6499__A1 _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7160__A2 _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5171__A1 _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7448__B1 _2692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7999__A1 _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6671__A1 _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5474__A2 _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5971_ _4362_ _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7710_ as2650.stack\[3\]\[5\] _2762_ _1045_ as2650.stack\[2\]\[5\] _2955_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4922_ _0293_ _0316_ _0365_ _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_8690_ net21 _3839_ _3867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_127_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8176__A1 _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7641_ _2886_ _2887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4853_ _0295_ _0296_ _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7923__A1 _2706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5908__I _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4812__I _4391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7572_ as2650.stack\[4\]\[2\] _2819_ _2694_ as2650.stack\[5\]\[2\] _2820_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4784_ _4363_ _4364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_18_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6523_ _4361_ _1845_ _1846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_140_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6454_ _1767_ _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7151__A2 _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4968__B _4146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7344__B _2599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5405_ as2650.r0\[1\] _0764_ _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5643__I _4063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6385_ _1632_ _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8124_ _0714_ _3263_ _3354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5336_ _4138_ _0738_ _0775_ _0006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8055_ _1381_ _3262_ _3288_ _1267_ _3289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_87_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5267_ _0328_ _0706_ _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7454__A3 _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7006_ as2650.addr_buff\[1\] _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_5_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5198_ _0638_ _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6414__A1 _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6414__B2 as2650.stack\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8957_ _0118_ clknet_leaf_56_wb_clk_i as2650.stack\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4976__A1 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7908_ as2650.pc\[11\] _0726_ _3147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8888_ _0049_ clknet_leaf_50_wb_clk_i as2650.stack\[1\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8167__A1 _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8622__C _3175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7839_ _2685_ _3080_ _2927_ _3081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7914__A1 _2796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6717__A2 _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7914__B2 _3152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4728__A1 _4289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7390__A2 _2580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6193__A3 _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5153__A1 _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5553__I _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8069__C _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4900__A1 _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8642__A2 _3819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6653__A1 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8085__B _3316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9039__CLK clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_75_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7905__A1 as2650.addr_buff\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5728__I _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4632__I _4212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5392__A1 as2650.r0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6987__C _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5144__A1 _4270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6892__A1 _1979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6170_ _1546_ _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5121_ as2650.r0\[2\] _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5447__A2 _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5052_ as2650.holding_reg\[4\] _0492_ _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_84_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6508__B _1830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8811_ _2307_ _2517_ _3978_ _3979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_77_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6947__A2 _2239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4958__A1 _4129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8742_ _1399_ _2550_ _2677_ _3915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_81_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5954_ _4087_ _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8149__A1 _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4905_ _0348_ _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8673_ _3852_ _1388_ _3853_ _3854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5885_ _0589_ _4308_ _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7624_ _2857_ _2859_ _2867_ _2870_ _2465_ _2871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4836_ _4415_ _4416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7372__A2 _2615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7555_ _0290_ _2803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5383__A1 _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4767_ _4343_ _4346_ _4347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6506_ _1809_ _1829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7486_ _1078_ _2735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8321__A1 net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7124__A2 _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4698_ _4278_ _4279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6437_ _1767_ _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6883__A1 as2650.r123_2\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6368_ _1714_ _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8107_ _2177_ _3245_ _3337_ _2730_ _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_130_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5319_ as2650.r0\[4\] _0464_ _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9087_ _0248_ clknet_leaf_26_wb_clk_i net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8624__A2 _3558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6299_ _1661_ _1662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6635__A1 _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5438__A2 _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8038_ _2898_ _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_103_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4717__I _4297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8388__A1 _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6938__A2 _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6932__I _2207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_45_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4949__A1 _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5610__A2 _4309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7363__A2 _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8560__A1 _3579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5992__B _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5374__A1 _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5126__A1 _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5283__I net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6874__A1 _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7418__A3 _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7003__I _2293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7051__A1 _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5601__A2 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_32_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5670_ _1094_ _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8551__A1 _3089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5365__A1 _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4621_ _4192_ _4077_ _4202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_124_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7340_ _2449_ _2596_ _2434_ _2542_ _2597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_11_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4552_ _4125_ _4127_ _4130_ _4132_ _4133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__8303__A1 _4090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7106__A2 _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6510__C _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6289__I _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7271_ _2530_ _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4483_ as2650.ins_reg\[5\] _4064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9010_ _0171_ clknet_leaf_80_wb_clk_i as2650.r123\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6865__A1 _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6222_ _1592_ _1160_ _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_49_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6153_ as2650.r123_2\[3\]\[2\] _1536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8606__A2 _3525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5104_ _0432_ _0537_ _0545_ _4204_ _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_83_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6084_ _4285_ _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4537__I _4033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7290__A1 _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5035_ _0474_ _0475_ _0477_ _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__8009__I _3243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5840__A2 _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6986_ _1057_ _2276_ _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__8790__A1 _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5937_ _0384_ _1320_ _0496_ _0497_ _1323_ _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_8725_ _4329_ _4354_ _3898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8656_ _3837_ _3840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5868_ _1262_ _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8542__A1 _3515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7345__A2 _2592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7607_ _2446_ _2834_ _2854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5356__A1 _4264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4819_ _4395_ _4398_ _4399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8587_ _1114_ _3480_ _3780_ _3498_ _3781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_107_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5799_ _1109_ _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7538_ as2650.pc\[2\] _0347_ _2786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_33_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7469_ _2708_ _2715_ _2718_ _2719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput13 net50 io_oeb[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_123_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput24 net24 io_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput35 net35 io_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_66_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7281__A1 _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7033__A1 _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8871__CLK clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8781__A1 _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5595__A1 as2650.r123\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8533__A1 _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6075__A2 _4108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5897__B _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6840_ _1386_ _1839_ _2155_ _1816_ _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_74_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6505__C _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6771_ _2075_ _2089_ _2090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5586__A1 as2650.stack\[7\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8510_ _3702_ _3706_ _3707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5722_ _1083_ _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8524__A1 _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7327__A2 _2574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8441_ _3639_ _0587_ _3640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5338__A1 _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5653_ _1051_ _1082_ _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4604_ _4147_ _4184_ _4185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8372_ _0348_ _0330_ _3573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5584_ _1014_ _1015_ _1016_ _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_102_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7323_ _2579_ _2564_ _2580_ _2581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4535_ _4043_ _4115_ _4075_ _4116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_117_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6838__A1 _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7254_ _2307_ _2513_ _2518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4466_ _4046_ _4047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_132_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6205_ _1575_ _1576_ _1579_ _0071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7185_ net25 _1553_ _2456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6136_ _1265_ _1517_ _1521_ _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7263__A1 _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6066__A2 _4116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6067_ _1450_ _1452_ _1453_ _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_3207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8894__CLK clknet_leaf_52_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5813__A2 _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5018_ _4139_ _0413_ _0460_ _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_96_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6482__I _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5577__A1 _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5098__I _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6969_ _1072_ _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8708_ _3880_ _3881_ _3882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8515__A1 _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8639_ _1205_ _3820_ _3826_ _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_139_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4552__A2 _4127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6829__A1 _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8358__B _3559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5501__A1 _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6057__A2 _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7254__A1 _2307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8805__C _2639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5804__A2 _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6392__I _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4905__I _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8754__A1 _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7557__A2 _4384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7309__A2 _2344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4791__A2 as2650.addr_buff\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4543__A2 _4123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8809__A2 _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input1_I io_in[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6048__A2 _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8990_ _0151_ clknet_leaf_68_wb_clk_i as2650.r123_2\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_68_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7941_ _2306_ _3178_ _3179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_83_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7872_ _3111_ _3084_ _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_51_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6823_ _0646_ _1819_ _2139_ _1815_ _2140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6220__A2 _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6754_ _2034_ _2047_ _2073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7347__B _2603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5705_ _0998_ _1099_ _1100_ _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_52_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6685_ _2003_ _2005_ _2006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_104_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8424_ net32 _3460_ _3623_ _3624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5636_ _1064_ _1065_ _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8355_ _1473_ _3532_ _3556_ _3294_ _3557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5567_ as2650.stack\[3\]\[12\] _0948_ _0949_ _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7306_ _2326_ _2564_ _2565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4518_ _4065_ _4041_ _4099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8286_ _3488_ _3489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5498_ _0886_ _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7484__A1 _1612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7237_ _2490_ _2504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4449_ _4029_ as2650.cycle\[2\] _4030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7168_ _1063_ _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6039__A2 _4291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6119_ _1501_ _1504_ _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_19_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7099_ _0462_ _2135_ _2360_ _0738_ _2372_ _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_74_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9072__CLK clknet_leaf_41_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4725__I _4189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7539__A2 _2786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5970__A1 _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7011__I1 _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4525__A2 _4101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8088__B _3242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7475__A1 _2701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5486__B1 _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7227__A1 _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7778__A2 _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5005__A3 _4388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8270__C _3473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7950__A2 _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5466__I _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6470_ _1793_ _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5421_ _4138_ _0818_ _0859_ _0007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4516__A2 _4096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7681__I _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8140_ _3368_ _0713_ _3244_ _3369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5352_ _4205_ _0681_ _0790_ _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7466__A1 _4125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8071_ _3303_ _3258_ _1385_ _3304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5283_ net2 _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7022_ _2306_ _2302_ _2308_ _0159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9095__CLK clknet_leaf_55_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7218__A1 _4094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8973_ _0134_ clknet_leaf_35_wb_clk_i as2650.stack\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6441__A2 _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8017__I _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7924_ _2813_ _3146_ _3162_ _3163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8718__A1 _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7855_ _2296_ _3095_ _3096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_51_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7856__I as2650.addr_buff\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6806_ _2111_ _2123_ _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7786_ _2704_ _3029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4998_ _4201_ _0440_ _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6737_ _1807_ _2056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5952__A1 _4396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4755__A2 _4298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6668_ _1987_ _1988_ _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8407_ _1409_ _0516_ _3606_ _3607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
X_5619_ _4141_ _0504_ _0872_ _0874_ _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_87_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6901__B1 _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6599_ _1848_ _1920_ _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8338_ _3502_ _3538_ _3539_ _3540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__8249__A3 _3450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7457__A1 _2539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8269_ _2267_ _2489_ _3473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6000__I _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7209__A1 _2455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output40_I net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6968__B1 _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5060__B _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8709__A1 _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4994__A2 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8090__C _3321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7932__A2 _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5943__A1 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5286__I _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7696__A1 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6499__A2 _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7448__A1 as2650.stack\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_57_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_57_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__7448__B2 as2650.stack\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7006__I as2650.addr_buff\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7999__A2 _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8546__B _2458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6671__A2 _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4682__A1 _4261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8955__CLK clknet_leaf_43_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7620__A1 _2862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5970_ _1351_ _1356_ _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4921_ _0292_ _0364_ _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7640_ _1687_ net9 _2886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6187__A1 _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4852_ as2650.holding_reg\[2\] _0294_ _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_61_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7923__A2 _3142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7571_ _1191_ _2819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4783_ _4048_ _4055_ _4363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6522_ _1056_ _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7687__A1 as2650.pc\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6453_ _1620_ _1774_ _1781_ _0117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5404_ _0665_ _0842_ _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7344__C _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6384_ as2650.stack\[3\]\[3\] _1715_ _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8123_ _2431_ _0607_ _3352_ _1473_ _3353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_126_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5335_ as2650.r123\[1\]\[6\] _4413_ _0774_ _4316_ _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_86_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8100__A2 _2923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8054_ _3282_ _3286_ _3287_ _3288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5266_ _0679_ _0705_ _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6111__A1 _1496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8651__A3 _3832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7005_ _2295_ _0155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5197_ _0396_ _0536_ _0637_ _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7611__A1 _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8956_ _0117_ clknet_leaf_56_wb_clk_i as2650.stack\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7907_ _3143_ _3145_ _3146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_70_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4976__A2 _4021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8887_ _0048_ clknet_leaf_51_wb_clk_i as2650.stack\[1\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6178__A1 _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7838_ _3053_ _3061_ _3079_ _2462_ _3080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_12_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9110__CLK clknet_leaf_9_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7914__A2 _3142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4728__A2 _4308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5925__A1 _4186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7769_ as2650.stack\[2\]\[7\] _3012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_71_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6193__A4 _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7678__A1 _2823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5153__A2 _4021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4900__A2 _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7850__A1 _3089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8978__CLK clknet_leaf_77_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6653__A2 _1973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8085__C _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6405__A2 _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4806__I3 as2650.r123_2\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7905__A2 _3097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5916__A1 as2650.stack\[0\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5392__A2 _4414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7669__A1 _2813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5931__A4 _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7164__C _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5144__A2 _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6341__A1 _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6892__A2 _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_39_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5120_ _4148_ _0561_ _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8094__A1 _3271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5051_ _0490_ _0492_ _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_97_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6508__C _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8810_ _1435_ _3974_ _3975_ _3977_ _3978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_81_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8741_ _1383_ _3262_ _1362_ _3914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5953_ _4223_ _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4958__A2 _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5080__A1 _4012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4904_ _0347_ _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8672_ _1628_ _3843_ _3853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5884_ _1278_ _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7623_ _1406_ _2868_ _2869_ _2870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4835_ _4414_ _4415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7554_ _2793_ _2795_ _2801_ _2427_ _2802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5383__A2 _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_78_wb_clk_i_I clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4766_ _4344_ _4345_ _4346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_140_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6505_ _4224_ _1819_ _1827_ _1815_ _1828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_88_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7485_ _2733_ _2734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4697_ _4265_ _4277_ _4278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7124__A3 _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6436_ _1082_ _1766_ _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6883__A2 _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6367_ _1713_ _0969_ _1605_ _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4894__A1 _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5318_ _0335_ _0367_ _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8085__A1 _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8106_ _3328_ _3336_ _3276_ _3337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_103_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9086_ _0247_ clknet_leaf_25_wb_clk_i net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6298_ _1660_ _1661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7832__A1 _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6485__I _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8037_ _3271_ _4272_ _3272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5249_ as2650.holding_reg\[6\] _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_5_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_2_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_57_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8388__A2 _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8939_ _0100_ clknet_leaf_37_wb_clk_i as2650.stack\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4949__A2 _4389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5071__A1 _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5829__I _4073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5610__A3 _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8560__A2 _3752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5992__C _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6571__A1 _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5564__I as2650.r123\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5126__A2 _4415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9006__CLK clknet_leaf_77_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4885__A1 _4270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8076__A1 _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7823__A1 _3064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7051__A2 _2332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8000__A1 _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4620_ _4199_ _4201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4551_ _4131_ _4059_ _4132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8303__A2 _3505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7270_ _4287_ _2530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4482_ _4062_ _4063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6221_ _1591_ _1592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4876__A1 _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6152_ _1535_ _0062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8067__A1 _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5103_ _0540_ _4245_ _4227_ _0544_ _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_97_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7814__A1 _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6083_ _1339_ _1361_ _1469_ _1470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_26_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5034_ _0371_ _0374_ _0476_ _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7290__A2 _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7578__B1 _2822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6985_ _2275_ _1253_ _2276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_41_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8790__A2 _3920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8724_ _4329_ _4353_ _4169_ _3896_ _3897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_81_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5936_ _1321_ _1322_ _0386_ _0298_ _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_80_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8655_ _3835_ _3839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5867_ _1215_ _1261_ _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8542__A2 _3736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7606_ _2301_ _2261_ _2606_ _2852_ _2853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_107_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5356__A2 _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4818_ _4265_ _4397_ _4398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8586_ _3779_ _3780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_124_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5798_ _1190_ _1197_ _1199_ _0044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__9029__CLK clknet_leaf_17_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7537_ _2783_ _2784_ _2785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_108_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4749_ _4328_ _4329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6305__A1 _1667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7468_ _1439_ _2708_ _2717_ _2718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xoutput14 net14 io_oeb[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput25 net25 io_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_6419_ _1624_ _1749_ _1752_ as2650.stack\[2\]\[2\] _1755_ _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_66_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput36 net36 io_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_7399_ _2494_ _2651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4867__A1 _4171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8058__A1 _2336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7805__A1 _2831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_9069_ _0230_ clknet_leaf_38_wb_clk_i as2650.stack\[7\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6148__C _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7281__A2 _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5292__A1 _4370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7569__B1 _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7033__A2 _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8781__A2 _2657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8533__A2 _3728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6847__A2 _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4858__A1 as2650.holding_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7014__I _2293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7024__A2 _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8221__A1 _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5469__I _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6770_ _2078_ _2088_ _2089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5586__A2 _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5721_ _1104_ _1143_ _1144_ _0022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_94_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8524__A2 _3326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8440_ _0603_ _3639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6535__A1 _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5652_ _4110_ _1081_ _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7732__B1 _2975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4603_ _4162_ _4165_ _4183_ _4184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8371_ _3571_ _3572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5583_ as2650.stack\[0\]\[13\] _0904_ _0918_ as2650.stack\[1\]\[13\] _1016_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_117_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7322_ _2273_ _2580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4534_ _4114_ _4115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6838__A2 _1855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4465_ as2650.cycle\[7\] _4046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7253_ _1481_ _2517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6204_ _1578_ _1565_ _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7184_ _2392_ _2448_ _2452_ _2454_ _2455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_131_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6135_ _1518_ _1519_ _1520_ _1244_ _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__4548__I _4115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6066_ _4310_ _4116_ _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8464__B _2980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5017_ _0442_ _0453_ _0459_ _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8212__A1 as2650.stack\[7\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5379__I _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8763__A2 _3924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6968_ _1258_ _2256_ _2258_ _1359_ _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8707_ _1283_ _2550_ _2677_ _3881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5919_ _1207_ _1302_ _1308_ _0056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_74_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6899_ _0677_ _1905_ _2193_ as2650.r123_2\[1\]\[5\] _2201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8515__A2 _3484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5329__A2 _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8638_ as2650.stack\[4\]\[11\] _3823_ _3826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6526__A1 _1842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8569_ _3472_ _2286_ _3763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8279__A1 _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6829__A2 _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8358__C _3485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5501__A2 _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8451__A1 _3537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5265__A1 _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8203__A1 _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5017__A1 _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8754__A2 _2325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5568__A2 _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6517__A1 _4045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7714__B1 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5740__A2 _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4569__S _4010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7172__C _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8690__A1 net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6048__A3 _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5256__A1 _4343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5256__B2 _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6583__I _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7940_ _3143_ _3145_ _3178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7871_ as2650.pc\[10\] _3111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_63_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5008__A1 _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5199__I _4193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6822_ _4223_ _1968_ _1818_ _2138_ _2139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7628__B _2791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6753_ _2049_ _2052_ _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5704_ _1129_ _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6508__A1 _4272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6684_ _1931_ _1958_ _2004_ _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8423_ _2459_ _3617_ _3622_ _3485_ _3623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_34_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5635_ as2650.addr_buff\[7\] _4124_ _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7181__A1 _2450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8354_ _3534_ _3536_ _3527_ _3537_ _3555_ _3556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_30_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5566_ _0517_ _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7305_ _2562_ _2563_ _2564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4517_ _4089_ _4092_ _4097_ _4098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_2_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8285_ _3459_ _3488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5497_ _0934_ _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8681__A1 _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7236_ _2500_ _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4448_ as2650.cycle\[3\] _4029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8861__CLK clknet_leaf_46_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7167_ _4194_ _2439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8433__A1 _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6118_ _1502_ _1387_ _4389_ _0348_ _1503_ _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7098_ as2650.r123\[2\]\[6\] _2364_ _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5247__A1 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6493__I _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6049_ _1341_ _4296_ _4331_ _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__5798__A2 _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8736__A2 _3906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6747__A1 _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7944__B1 _3181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5837__I _4214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4741__I _4321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5970__A2 _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8369__B _3464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4525__A3 _4105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4930__B1 _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8672__A1 _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8424__A1 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7227__A2 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5238__A1 _4138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5789__A2 _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6738__A1 _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5005__A4 _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5747__I _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5410__A1 _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7163__A1 net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5420_ as2650.r123\[1\]\[7\] _4304_ _0858_ _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_127_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8884__CLK clknet_leaf_52_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6910__A1 _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5351_ _4228_ _0782_ _0789_ _4205_ _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5482__I _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8070_ _1365_ _3303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5282_ _4247_ _0721_ _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_88_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7466__A2 _4151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7021_ _2307_ _2304_ _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8415__A1 _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7218__A2 _2485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8972_ _0133_ clknet_leaf_35_wb_clk_i as2650.stack\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7202__I _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout52_I net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7923_ _2706_ _3142_ _3154_ _3160_ _3161_ _3162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__6441__A3 _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8718__A2 _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7854_ _3063_ _3065_ _3095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6729__A1 _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8461__C _3659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7926__B1 _3163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7358__B _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6805_ _2118_ _2122_ _2123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7785_ _2576_ _3025_ _3027_ _3028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5657__I _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5401__A1 _4148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4997_ _4205_ _4390_ _0439_ _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4561__I _4141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8033__I _2547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6736_ _1962_ _2026_ _2027_ _2055_ _0126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7154__A1 _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6667_ _0337_ _1936_ _0470_ _4209_ _1988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_104_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8406_ _3604_ _3605_ _3606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5618_ _1047_ _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5165__B1 _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6598_ _4359_ _1907_ _1916_ _1919_ _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_121_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8337_ _4392_ _4358_ _3539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5549_ _0946_ _0983_ _0984_ _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8103__B1 _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7457__A2 _2706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8268_ _2272_ _3472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5468__A1 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7219_ _4057_ _2484_ _2487_ _2479_ _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_63_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8199_ _1599_ _3416_ _3417_ _3418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4736__I _4316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8208__I _3411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6968__A1 _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6968__B2 _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output33_I net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8709__A2 _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5640__A1 _4170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5995__C _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7393__A1 _2430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7696__A2 _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_29_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8645__A1 _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_3_6_0_wb_clk_i clknet_0_wb_clk_i clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_69_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_0_wb_clk_i_I wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4646__I _4226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_26_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_26_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_77_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6959__A1 _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8562__B _3098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6861__I _2165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4920_ _0317_ _0327_ _0363_ _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4851_ as2650.holding_reg\[2\] _0294_ _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6187__A2 _1563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5477__I _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7570_ as2650.stack\[7\]\[2\] _2762_ _1046_ as2650.stack\[6\]\[2\] _2818_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4782_ _4361_ _4362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5934__A2 _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_68_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7906__B _3144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6521_ _0864_ _1843_ _1805_ _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_53_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7687__A2 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7625__C _2537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6452_ as2650.stack\[1\]\[2\] _1768_ _1780_ _1773_ _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__5698__A1 as2650.r123\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5403_ _0524_ _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__9062__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6383_ _1628_ _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8122_ _1287_ _1363_ _3350_ _3351_ _2724_ _3352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_142_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5334_ _0773_ _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_115_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8053_ _4417_ _0934_ _4078_ _3287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5265_ _0582_ _0583_ _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6111__A2 _4249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7004_ _2252_ _1559_ _2294_ _2295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5196_ _0636_ _4295_ _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4673__A2 _4239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5870__A1 _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8028__I _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7611__A2 _1612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8955_ _0116_ clknet_leaf_43_wb_clk_i as2650.stack\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8472__B _3468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7906_ _3064_ _3034_ _3144_ _2545_ _3145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_71_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8886_ _0047_ clknet_leaf_52_wb_clk_i as2650.stack\[1\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7837_ _0925_ _2961_ _3060_ _3077_ _3078_ _3079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__6178__A2 _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7768_ _1655_ _3010_ _3011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5925__A2 _4355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6719_ _1993_ _1994_ _2039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7699_ _2851_ _2943_ _2944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7678__A2 _2923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5689__A1 as2650.r123\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6011__I _4243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8627__A1 _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7551__B _1440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5850__I _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7602__A2 _2848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6405__A3 _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8563__B1 _3757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5916__A2 _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9085__CLK clknet_leaf_24_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7118__A1 _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7669__A2 _2906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5246__B _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8618__A1 _3173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6856__I _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8094__A2 _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5050_ _0491_ _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5852__A1 _4032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4655__A2 _4235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8292__B _2750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5604__A1 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8740_ _3303_ _0717_ _2492_ _3912_ _3313_ _3913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_81_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5952_ _4396_ _1311_ _1314_ _1338_ _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_92_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4903_ net7 _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
X_8671_ _3837_ _3852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5883_ _1225_ _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7622_ _2745_ _2869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4834_ as2650.r123\[0\]\[1\] as2650.r123_2\[0\]\[1\] _4008_ _4414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5000__I _4270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7553_ _2797_ _2799_ _2800_ _2801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_53_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7109__A1 _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4765_ _4177_ _4158_ _4162_ _4345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__6580__A2 _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6504_ _4239_ _1821_ _1826_ _1818_ _1827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7355__C _2334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4591__A1 _4141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7484_ _1612_ _1666_ _2733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4696_ _4275_ _4276_ _4277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6435_ _1043_ _1194_ _1766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_128_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5540__B1 _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6366_ _0910_ _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_66_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4995__B _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7371__B _2626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8105_ _1569_ _0543_ _2651_ _0428_ _3335_ _3336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_143_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5317_ _0417_ _0369_ _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9085_ _0246_ clknet_leaf_24_wb_clk_i net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5670__I _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8085__A2 _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6297_ _1592_ _1147_ _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6096__A1 _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8036_ _2626_ _3271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7832__A2 _3058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5248_ _0682_ _0687_ _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_76_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5843__A1 _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5179_ _0317_ _0619_ _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_84_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8388__A3 _2569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8938_ _0099_ clknet_leaf_42_wb_clk_i as2650.stack\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_43_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5071__A2 _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7348__A1 _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8869_ _0030_ clknet_leaf_49_wb_clk_i as2650.stack\[6\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5610__A4 _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6006__I _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6571__A2 _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8945__CLK clknet_leaf_56_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7520__A1 _2760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4885__A2 _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8076__A2 _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5834__A1 _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7587__A1 _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7300__I _2409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7339__A1 _2594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8000__A2 _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4550_ _4022_ _4131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4481_ as2650.ins_reg\[2\] _4062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7511__A1 _2724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6220_ _0861_ _1093_ _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_83_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6586__I _1842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4876__A2 _4388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6151_ as2650.r123_2\[3\]\[1\] _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8067__A2 _2822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_41_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_41_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6078__A1 _4037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5102_ _4245_ _0543_ _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6082_ _1415_ _1468_ _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5825__A1 _4006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5033_ _0333_ _0373_ _4320_ _0372_ _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7578__A1 _2790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7578__B2 _2823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8306__I _3468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6984_ _4053_ _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_65_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8723_ _0486_ _4184_ _3895_ _3896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5935_ _4156_ _4169_ _4344_ _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8750__B _2335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8654_ _3837_ _3838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5866_ _1049_ _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6002__A1 _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7605_ _1406_ _2851_ _2852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4817_ as2650.ins_reg\[4\] _4396_ _4397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8585_ _3040_ _3125_ _3493_ _3778_ _3779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_33_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7750__A1 _2857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5797_ as2650.stack\[1\]\[8\] _1198_ _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8968__CLK clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7536_ _2711_ _2748_ _2784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4748_ _4114_ _4238_ _4327_ _4328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7467_ _4242_ _2716_ _2717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7502__A1 as2650.addr_buff\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4679_ _4088_ _4260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6418_ _1744_ _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput15 net15 io_oeb[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_116_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput26 net26 io_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_7398_ _2640_ _2650_ _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xoutput37 net37 io_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_118_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4867__A2 _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8058__A2 _4400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6349_ _1702_ _0092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6069__A1 _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6069__B2 _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9068_ _0229_ clknet_leaf_42_wb_clk_i as2650.stack\[7\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8019_ _0905_ _3252_ _3253_ _3254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_76_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5292__A2 _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7569__A1 as2650.stack\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7569__B2 as2650.stack\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4744__I _4137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7741__A1 _1650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4555__A1 _4024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8835__B _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8221__A2 _3412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6232__A1 _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_51_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7980__A1 _2701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5720_ as2650.stack\[3\]\[14\] _1086_ _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5651_ _1067_ _1068_ _1071_ _1080_ _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_104_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5485__I _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6535__A2 _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7732__A1 _2885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7732__B2 _2892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4602_ _4168_ _4169_ _4165_ _4182_ _4183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_8370_ _4097_ _3571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5582_ as2650.stack\[2\]\[13\] _0969_ _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7321_ _2574_ _2579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_102_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4533_ _4113_ _4114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7252_ _2516_ _0181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4464_ _4027_ _4038_ _4044_ _4045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_116_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6203_ _1577_ _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7183_ _4301_ _4084_ _1079_ _2453_ _2398_ _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_113_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6134_ _1076_ _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7799__A1 _2892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6065_ _1451_ _4193_ _1436_ _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6471__A1 _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5016_ _0317_ _0458_ _0292_ _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8036__I _2626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6967_ _1352_ _2257_ _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5918_ as2650.stack\[0\]\[12\] _1304_ _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8706_ _3873_ _3877_ _3879_ _3880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6898_ _2068_ _2192_ _2200_ _0143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8637_ _1203_ _3820_ _3825_ _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5849_ _1240_ _1242_ _1243_ _0350_ _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__7723__A1 _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6526__A2 _1824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8568_ _3595_ _3762_ _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7519_ _2316_ _2767_ _2768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8279__A2 _2571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8499_ _3603_ _3695_ _3696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4739__I _4319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7115__I _4250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8451__A2 _3631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5265__A2 _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8754__A3 _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7962__A1 _2599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6517__A2 _4061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7714__A1 as2650.stack\[7\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4649__I _4229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5254__B _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8690__A2 _3839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8442__A2 _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6453__A1 _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6085__B _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7870_ _1114_ _2775_ _3110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5008__A2 _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6205__A1 _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6821_ _1373_ _1823_ _2137_ _1836_ _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_36_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6752_ _1801_ _2071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4767__A1 _4343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5703_ _1128_ _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6683_ _1933_ _1957_ _2004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7705__A1 _1440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6508__A2 _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8422_ _1639_ _3558_ _3621_ _3622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4519__A1 _4062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5634_ _1056_ _1063_ _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5716__B1 _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8353_ _3472_ _3554_ _3555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5565_ _0998_ _0942_ _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7304_ _4194_ _4056_ _2563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7363__C _2618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4516_ _4093_ _4096_ _4097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8284_ _3338_ _3487_ _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8130__A1 _3324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5496_ _0926_ _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7235_ _2502_ _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4447_ as2650.cycle\[7\] as2650.cycle\[6\] as2650.cycle\[5\] as2650.cycle\[4\] _4028_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_132_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7166_ _2437_ _2438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6117_ _0540_ _0427_ _0601_ _1372_ _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7097_ _0651_ _2360_ _2371_ _0171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6048_ _4007_ _1284_ _1217_ _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_3017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7819__B _2770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7999_ _1443_ _2562_ _1343_ _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7944__A1 _2796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6747__A2 _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7944__B2 _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4758__A1 _4156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6014__I _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5183__A1 as2650.holding_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4930__A1 _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8121__A1 _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5486__A2 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8424__A2 _3460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7227__A3 _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5238__A2 _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5521__C _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6986__A2 _2276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8188__A1 _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_58_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8360__A1 _3338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7163__A2 _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6910__A2 _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7183__C _2398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4921__A1 _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5350_ _0785_ _4246_ _4228_ _0788_ _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__8112__A1 _2623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5281_ _0601_ _0720_ _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_82_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7020_ _1410_ _2307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6426__A1 _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6426__B2 as2650.stack\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8971_ _0132_ clknet_leaf_35_wb_clk_i as2650.stack\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7922_ _2472_ _3150_ _3157_ _2647_ _2537_ _3161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_36_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8179__A1 _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7853_ _2782_ _3087_ _3093_ _2789_ _3094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_110_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7926__A1 _2894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8314__I _2409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6804_ _2120_ _2121_ _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7784_ _2558_ _2804_ _1430_ _2312_ _3026_ _3027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4996_ _4228_ _0428_ _0438_ _4380_ _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_51_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6735_ _1867_ _2054_ _2055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5952__A3 _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6666_ _0756_ _1986_ _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7154__A2 _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8351__A1 _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7374__B _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8405_ _2899_ _0457_ _3540_ _3541_ _3566_ _3605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_104_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5617_ _1046_ _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5165__A1 _4077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5673__I _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6597_ _4374_ _1918_ _1906_ _1919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_30_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8336_ _4391_ _4358_ _3538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5548_ _0366_ _0870_ _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_3_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8103__A1 _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_opt_3_0_wb_clk_i clknet_3_6_0_wb_clk_i clknet_opt_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_117_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8103__B2 _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8267_ _3464_ _3467_ _3470_ _2256_ _3471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_65_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5479_ as2650.stack\[0\]\[8\] _0904_ _0908_ as2650.stack\[1\]\[8\] _0916_ _0917_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_133_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6665__A1 _4208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5468__A2 _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7218_ _4094_ _2485_ _2484_ _2487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8198_ _3408_ _3417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7149_ _1451_ _1423_ _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6417__A1 _1611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6968__A2 _2256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7090__A1 _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6009__I _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5640__A2 _4044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output26_I net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5848__I _4027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8590__A1 net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7393__A2 _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xfanout50 net13 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_23_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7145__A2 _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8099__C _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8645__A2 _3821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6656__A1 _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5532__B _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6959__A2 _2207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_66_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_66_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_92_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4662__I _4242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8030__B1 _3264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4850_ _4388_ _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8851__CLK clknet_leaf_66_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4781_ _4088_ _4361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6520_ _0865_ _1843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6451_ _1623_ _1750_ _1766_ _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_70_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5402_ _0837_ _0838_ _0840_ _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_31_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9170_ net47 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6382_ _1675_ _1722_ _1725_ _1726_ _0101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_86_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8121_ _1479_ _1386_ _4101_ _3351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5333_ _0741_ _0772_ _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__8636__A2 _3823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8737__C _3869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8052_ _0887_ _2767_ _3285_ _3286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5264_ _0599_ _0703_ _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_69_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7003_ _2293_ _2294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__4837__I _4416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5195_ as2650.holding_reg\[5\] _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5870__A2 _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7611__A3 _2703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8954_ _0115_ clknet_leaf_47_wb_clk_i as2650.stack\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7905_ as2650.addr_buff\[0\] _3097_ as2650.addr_buff\[2\] _3144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8885_ _0046_ clknet_leaf_52_wb_clk_i as2650.stack\[1\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5668__I _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4572__I _4152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7836_ _2824_ _3053_ _3078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6178__A3 _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8572__A1 _3731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7375__A2 _2628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7767_ as2650.pc\[6\] as2650.pc\[5\] _2930_ _3010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4979_ as2650.r123\[1\]\[4\] as2650.r123\[0\]\[4\] as2650.r123_2\[1\]\[4\] as2650.r123_2\[0\]\[4\]
+ _4002_ _0339_ _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__5925__A3 _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6718_ _1949_ _2037_ _2038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_71_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8324__A1 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7127__A2 _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7698_ _2940_ _2904_ _2941_ _2943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_71_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5138__A1 _4324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6649_ _1495_ _1837_ _1909_ _1969_ _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_118_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8319_ _1615_ _3490_ _3521_ _2572_ _3522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_65_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7551__C _2798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8874__CLK clknet_leaf_46_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4482__I _4062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8563__A1 _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8563__B2 _3654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7118__A2 _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5129__A1 _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6877__A1 _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6202__I _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5246__C _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8838__B _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7234__S _2501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5301__A1 _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5852__A2 _4118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5065__B1 _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5951_ _1316_ _1319_ _1337_ _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_94_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4902_ _0345_ _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8670_ _3835_ _3851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5882_ _1228_ _1239_ _1250_ _1276_ _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__7357__A2 _4121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8554__A1 _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7621_ _2809_ _2868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4833_ _4303_ _4413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7552_ _1052_ _2787_ _2800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4764_ _4333_ _4336_ _4344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__7109__A2 _4170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6580__A3 _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6503_ _4243_ _1823_ _1825_ _1820_ _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_119_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4591__A2 _4171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7483_ _2461_ _2732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4695_ _4057_ as2650.idx_ctrl\[0\] _4276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6434_ _1667_ _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6365_ _1711_ _1712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8104_ _1411_ _1395_ _3333_ _3334_ _2586_ _3335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_118_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5316_ _0336_ _0467_ _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9084_ _0245_ clknet_leaf_25_wb_clk_i net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6296_ _1654_ _1637_ _1659_ _0082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5172__B _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8035_ _3269_ _3270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4567__I as2650.r0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6096__A2 _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7293__A1 _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5247_ _0624_ _0686_ _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5843__A2 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5178_ _0618_ _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7045__A1 _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8793__A1 _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8937_ _0098_ clknet_leaf_61_wb_clk_i as2650.r123\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4654__I0 as2650.r123\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8868_ _0029_ clknet_leaf_46_wb_clk_i as2650.stack\[5\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7348__A2 _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7819_ _2780_ _3060_ _2770_ _3061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_24_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8799_ _1859_ _1220_ _3967_ _3968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_71_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6859__A1 _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6022__I _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6859__B2 as2650.stack\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8658__B _3839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7520__A2 _2734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5861__I _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8377__C _2622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7284__A1 _2434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8393__B _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7587__A2 _2833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8784__A1 _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5598__A1 as2650.stack\[7\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9052__CLK clknet_leaf_66_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8536__A1 _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7339__A2 _2595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7028__I _2311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4480_ _4048_ _4049_ _4056_ _4060_ _4061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_116_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7511__A2 _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5771__I _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6150_ _1534_ _0061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6078__A2 _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5101_ _0492_ _0542_ _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_83_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6081_ _1432_ _1448_ _1456_ _1467_ _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5032_ _0469_ _0471_ _0472_ _0473_ _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5825__A2 _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_81_wb_clk_i clknet_3_0_0_wb_clk_i clknet_leaf_81_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_66_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_10_wb_clk_i clknet_3_2_0_wb_clk_i clknet_leaf_10_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_93_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7578__A2 _2815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6983_ _2268_ _2273_ _1449_ _4284_ _2274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_94_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8722_ _4325_ _4159_ _3895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5934_ _4329_ _0305_ _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8527__A1 _3051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5865_ _1259_ _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8653_ _0864_ _3837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6002__A2 _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4850__I _4388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7604_ _2260_ _2851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4816_ as2650.ins_reg\[5\] as2650.ins_reg\[6\] as2650.ins_reg\[7\] _4396_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__and3_1
X_8584_ _3126_ _3777_ _3778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5796_ _1196_ _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7750__A2 _2985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7535_ as2650.pc\[1\] net6 _2783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5761__A1 _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4747_ _4326_ _4113_ _4327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7466_ _4125_ _4151_ _2716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4678_ _4189_ _4200_ _4256_ _4258_ _4259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__7502__A2 _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6417_ _1611_ _1746_ _1754_ _0108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8909__D _0070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7397_ _2531_ _2408_ _2649_ _2650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5681__I _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput16 net16 io_oeb[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_89_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput27 net27 io_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_122_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput38 net38 io_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_122_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6348_ as2650.r123\[3\]\[1\] _1702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6069__A2 _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6069__B3 _4196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9067_ _0228_ clknet_leaf_38_wb_clk_i as2650.stack\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6279_ _1644_ _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5816__A2 _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8018_ _0887_ _3253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7018__A1 _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9075__CLK clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5029__B1 _4416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8766__A1 _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6017__I _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8518__A1 net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5856__I as2650.halted vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8912__CLK clknet_leaf_9_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5752__A1 as2650.stack\[6\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5807__A2 _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8757__A1 _4308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4491__A1 _4063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6232__A2 _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4871__S _4146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8509__A1 _3602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5991__A1 _4007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5650_ _4142_ _1072_ _1079_ _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7732__A2 _2968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4601_ _4171_ _4156_ _4172_ _4176_ _4181_ _4182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5581_ as2650.stack\[3\]\[13\] _0948_ _0950_ _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7320_ _2573_ _2575_ _2577_ _2578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4532_ _4062_ as2650.ins_reg\[3\] _4113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_8_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7496__A1 _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7251_ _0395_ _2515_ _2501_ _2516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_89_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4463_ _4040_ _4043_ _4044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6202_ _1224_ _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7182_ _4054_ _4122_ _2453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_28_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9098__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6133_ _1488_ _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7799__A2 _3024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6064_ _4083_ _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5015_ _0457_ _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6471__A2 _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8935__CLK clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6966_ _1241_ _1078_ _2257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7377__B _2590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8705_ _4207_ _1859_ _1220_ _2280_ _3878_ _3879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5917_ _1205_ _1301_ _1307_ _0055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5982__A1 _4164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6897_ as2650.r123_2\[1\]\[4\] _2189_ _2199_ _2200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_70_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8636_ as2650.stack\[4\]\[10\] _3823_ _3825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5848_ _4027_ _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_107_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8567_ net51 _3460_ _3761_ _3762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5779_ _1118_ _1180_ _1185_ _0039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_120_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7518_ _2761_ _2763_ _2766_ _2767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8498_ _1519_ _0797_ _3694_ _3695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_108_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7449_ as2650.stack\[0\]\[0\] _1194_ _2695_ as2650.stack\[1\]\[0\] _0923_ _2699_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_107_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9119_ _0280_ clknet_leaf_45_wb_clk_i as2650.psl\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8227__I _3436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8739__A1 _3911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6970__I _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7411__A1 _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7411__B2 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7962__A2 _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_48_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7478__A1 _2438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7750__B _2993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8958__CLK clknet_leaf_47_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6453__A2 _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4464__A1 _4027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7402__A1 _4048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6205__A2 _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6820_ _2136_ _1853_ _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6751_ as2650.r123_2\[2\]\[4\] _2069_ _2070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5964__A1 _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5496__I _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5702_ as2650.pc\[12\] _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6682_ _1999_ _2002_ _2003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__7705__A2 _2948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8421_ _1689_ _3525_ _3620_ _2473_ _2687_ _3621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_104_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5633_ _1057_ _1062_ _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5716__A1 as2650.pc\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4519__A2 _4099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5716__B2 as2650.r123_2\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8352_ _3546_ _3547_ _3553_ _3554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5564_ as2650.r123\[0\]\[4\] _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5192__A2 _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7303_ _2311_ _2561_ _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4515_ _4094_ _4095_ _4096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7469__A1 _2708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8283_ _3447_ _3460_ _3486_ _3487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5495_ as2650.r123\[0\]\[0\] _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8130__A2 _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7234_ as2650.holding_reg\[0\] _2492_ _2501_ _2502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4446_ _4026_ _4027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7165_ _1358_ _2323_ _2437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6116_ net6 _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_113_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7096_ _0288_ _2124_ _2368_ as2650.r123\[2\]\[5\] _2371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6047_ _1433_ _1394_ _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8047__I _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4455__A1 _4032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8491__B _3687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5400__S _4009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7998_ _4364_ _4060_ _1431_ _3232_ _2268_ _3233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_54_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9113__CLK clknet_leaf_43_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7944__A2 _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4758__A2 _4157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6949_ _2106_ _2229_ _2243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_74_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8619_ _3626_ _3810_ _3811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_127_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5183__A2 _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6380__A1 as2650.stack\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8121__A2 _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6965__I _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6683__A2 _1957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7632__A1 _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6435__A2 _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4997__A2 _4390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7796__I _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_4_wb_clk_i_I clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6199__A1 _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7935__A2 _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5946__A1 as2650.psl\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7699__A1 _2851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7163__A3 _2434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8112__A2 _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5280_ _0718_ _0719_ _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6123__A1 as2650.psl\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5712__C _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7623__A1 _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8970_ _0131_ clknet_leaf_34_wb_clk_i as2650.stack\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7921_ _2280_ _3159_ _2735_ _3160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_48_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7852_ _2788_ _3092_ _3093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_63_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7926__A2 _3142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6803_ _2073_ _2074_ _2089_ _2121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7783_ _2599_ _3011_ _2489_ _3026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5937__B2 _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4995_ _0431_ _4246_ _0432_ _0437_ _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6734_ _2028_ _2031_ _2053_ _2054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_108_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6665_ _4208_ _1935_ _1986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7154__A3 _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8404_ _0430_ _0457_ _3604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7374__C _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5616_ _1045_ _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5165__A2 _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6596_ _1917_ _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8335_ _3505_ _3537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5547_ _0966_ _0980_ _0982_ _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8103__A2 _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8266_ _1496_ _3469_ _3470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5478_ _0915_ _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7217_ _4058_ _2484_ _2486_ _2479_ _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__7862__A1 _2793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6665__A2 _1935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4429_ _4009_ _4010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8197_ _3415_ _3416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4676__A1 _4024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7148_ _4362_ _2416_ _2419_ _2420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_63_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7079_ _0868_ _1520_ _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_100_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7090__A2 _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5640__A3 _4214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7917__A2 _3155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5928__A1 _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6025__I _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xfanout51 net37 net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_126_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4600__A1 _4177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5864__I _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5400__I0 as2650.r123\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7853__A1 _2782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7605__A1 _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5092__A1 _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7908__A2 _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8030__A1 _3262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8030__B2 _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4780_ _4280_ _4359_ _4360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6592__A1 _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_35_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_35_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_144_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8333__A2 _2786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6450_ _1779_ _0116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6344__A1 _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5401_ _4148_ _0839_ _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6895__A2 _2192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6381_ _1679_ _1718_ _1719_ _1726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_114_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5332_ _0744_ _0771_ _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8120_ _3344_ _3349_ _3281_ _3350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_138_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7922__C _2537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7844__A1 _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8051_ _1511_ _3283_ _3284_ _0886_ _3285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5263_ _0615_ _0580_ _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_130_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7002_ _2254_ _2259_ _2279_ _2292_ _2293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_114_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5194_ _0627_ _0633_ _0634_ _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8953_ _0114_ clknet_leaf_59_wb_clk_i as2650.stack\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5949__I _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7904_ as2650.addr_buff\[3\] _3143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8884_ _0045_ clknet_leaf_52_wb_clk_i as2650.stack\[1\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7835_ _2592_ _3076_ _3077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7766_ _1657_ _2775_ _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4978_ _4213_ _0420_ _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5925__A4 _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6717_ _0533_ _2036_ _2037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7697_ _2940_ _2904_ _2941_ _2942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__8324__A2 net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5138__A2 _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6648_ _0357_ _1855_ _1967_ _1968_ _1969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_109_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6579_ _1875_ _1901_ _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_124_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4897__A1 _4213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8088__A1 _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8318_ _1360_ _3499_ _3520_ _3521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7832__C _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7835__A1 _2592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8249_ _2375_ _2666_ _3450_ _3452_ _3453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_121_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4821__A1 _4244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8012__A1 _4004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8563__A2 _3525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5377__A2 _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7771__B1 _2956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7295__B _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8315__A2 _3494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5129__A2 _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7826__A1 _1656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7314__I _2571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8251__A1 _2311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5065__A1 _4168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5065__B2 _4299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5950_ _1332_ _1333_ _1336_ _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8003__A1 _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4901_ _0344_ _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5881_ _1252_ _1257_ _1264_ _1275_ _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA__7357__A3 _4103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7620_ _2862_ _2865_ _2866_ _2867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4832_ _4139_ _4355_ _4411_ _4412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_107_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6565__A1 _4229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7551_ _1575_ _2593_ _1440_ _2798_ _2799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_53_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4763_ _4065_ _4298_ _4343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_144_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7109__A3 _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6502_ _4250_ _1824_ _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6317__A1 as2650.stack\[4\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4694_ as2650.idx_ctrl\[1\] _4058_ _4275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7482_ _2727_ _2731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6433_ _1654_ _1758_ _1764_ _0114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5009__I _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4879__A1 _4232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6364_ _1710_ _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5540__A2 _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7817__A1 _2891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8103_ _1381_ _1495_ _0714_ _3281_ _1395_ _3334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_142_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5315_ _0753_ _0754_ _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_66_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9083_ _0244_ clknet_leaf_24_wb_clk_i net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6295_ _1657_ _1604_ _1608_ _1658_ _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8034_ _1426_ _3269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8490__A1 _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6096__A3 _4128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7293__A2 _2550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5246_ _0494_ _0502_ _0623_ _0493_ _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_29_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5177_ _0512_ _0581_ _0584_ _0455_ _0617_ _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_68_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7045__A2 _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8242__A1 _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5056__B2 _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8793__A2 _3940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8936_ _0097_ clknet_leaf_71_wb_clk_i as2650.r123\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4803__A1 _4382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4654__I1 as2650.r123\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8867_ _0028_ clknet_leaf_49_wb_clk_i as2650.stack\[5\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8545__A2 _3739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7818_ _2781_ _3053_ _3059_ _2789_ _3060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_40_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5359__A2 _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7753__B1 _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8798_ _1405_ _2677_ _3967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7749_ _1412_ _2868_ _2990_ _2992_ _2869_ _2993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_61_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8004__B _3238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8481__A1 _3603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7284__A2 _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8841__CLK clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5589__I _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5047__A1 _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8784__A2 _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8991__CLK clknet_leaf_68_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5598__A2 _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8536__A2 _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5100_ _0433_ _0345_ _0444_ _0541_ _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8472__A1 _3667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6080_ _1457_ _1458_ _1461_ _1466_ _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_98_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5031_ _0469_ _0471_ _0472_ _0473_ _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5499__I _4108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8775__A2 _3938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6982_ _2269_ _2272_ _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8721_ _0315_ _3893_ _3894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5933_ _0388_ _0303_ _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_50_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_59_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8652_ _3835_ _3836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7647__C _2758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5864_ _1219_ _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7603_ _2843_ _2849_ _2850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6002__A3 _4390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4815_ _4394_ _4249_ _4395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8583_ _2546_ _3770_ _3777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5795_ _1196_ _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7534_ _2781_ _2782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4746_ as2650.holding_reg\[1\] _4326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5761__A2 _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8759__B _2467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7465_ _1597_ _2445_ _2709_ _2714_ _2715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_119_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4677_ _4257_ _4258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6416_ _1670_ _1749_ _1752_ as2650.stack\[2\]\[1\] _1745_ _1754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__8864__CLK clknet_leaf_53_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7396_ _2531_ _2411_ _2645_ _2648_ _2649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
Xoutput17 net17 io_oeb[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput28 net28 io_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_66_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput39 net39 io_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_118_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6347_ _1701_ _0091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8463__A1 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6069__A3 _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9066_ _0227_ clknet_leaf_42_wb_clk_i as2650.stack\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6278_ _1643_ _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8017_ _3251_ _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5229_ _0669_ _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7018__A2 _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8215__A1 as2650.stack\[7\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5029__A1 _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8766__A2 _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6777__A1 _1962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8919_ _0080_ clknet_leaf_33_wb_clk_i as2650.stack\[5\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_38_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5201__A1 _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5752__A2 _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6701__A1 _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8454__A1 _2949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5268__A1 _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5268__B2 _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_77_wb_clk_i_I clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8206__A1 _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8757__A2 _3928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8509__A2 _3705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5991__A2 _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4600_ _4177_ _4159_ _4180_ _4181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8887__CLK clknet_leaf_51_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5743__A2 _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5580_ as2650.r123\[0\]\[5\] _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6940__A1 _2023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4531_ _4110_ _4111_ _4112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7496__A2 _2708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7250_ _1627_ _2513_ _2514_ _2515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_89_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8693__A1 _2431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4462_ _4042_ _4043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6201_ _1565_ _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7181_ _2450_ _2451_ _2452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6132_ as2650.psl\[7\] _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5259__A1 _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6063_ _1342_ _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5014_ _0454_ _0400_ _0446_ _0455_ _0456_ _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_113_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6759__A1 _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7420__A2 _2669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6965_ _2255_ _2256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_54_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5431__A1 _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5957__I _4143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8704_ _1457_ _1458_ _3878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5916_ as2650.stack\[0\]\[11\] _1304_ _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7971__A3 _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6896_ _0577_ _2012_ _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_62_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6281__C _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5982__A2 _4099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8635_ _1200_ _3820_ _3824_ _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7184__A1 _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5847_ _1241_ _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6526__A4 _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8566_ _3756_ _3760_ _3488_ _3761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5734__A2 _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6931__A1 as2650.r123_2\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5778_ as2650.stack\[2\]\[10\] _1183_ _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7517_ as2650.stack\[2\]\[1\] _2691_ _2765_ _0922_ _2766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4729_ _4231_ _4310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__9164__I net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8497_ _3673_ _3676_ _3693_ _3694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8684__A1 _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7448_ as2650.stack\[3\]\[0\] _2697_ _2692_ as2650.stack\[2\]\[0\] _2698_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_68_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9042__CLK clknet_leaf_29_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7379_ _1252_ _2613_ _2634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_81_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8436__A1 _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9118_ _0279_ clknet_leaf_46_wb_clk_i as2650.psl\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9049_ _0210_ clknet_leaf_40_wb_clk_i as2650.pc\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6998__A1 _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6456__C _1773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4473__A2 _4033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8739__A2 _2488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7411__A2 _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8243__I net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5725__A2 _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6922__A1 _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8675__A1 _3851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7750__C _2592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7322__I _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4464__A2 _4038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6750_ _1864_ _2069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5964__A2 _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5701_ _1087_ _1126_ _1127_ _0019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6681_ _2000_ _2001_ _2002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8420_ _2884_ _2890_ _3619_ _3620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7705__A3 _2949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5632_ _1058_ _4121_ _4119_ _1061_ _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__5177__B1 _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6913__A1 _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7925__C _2687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8351_ _1404_ _3509_ _3552_ _2625_ _3553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__9065__CLK clknet_leaf_40_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5563_ _0997_ _0011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7302_ _4090_ _4056_ _2561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6401__I _1656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4514_ as2650.addr_buff\[5\] _4095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7469__A2 _2715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8666__A1 _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8282_ _3461_ _3482_ _3484_ _1765_ _3485_ _3486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5494_ _4283_ _0871_ _0878_ _0931_ _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_117_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7233_ _2500_ _2501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4445_ _4025_ _4026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8418__A1 _2851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7164_ _2429_ _2432_ _2435_ _1362_ _2436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_67_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6115_ _1499_ _0716_ _1482_ _1500_ _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_99_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7095_ _0558_ _2360_ _2370_ _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6046_ _4084_ _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4455__A2 _4035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5652__A1 _4110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6995__A4 _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7997_ _2860_ _4396_ _1843_ _4096_ _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6948_ as2650.r123_2\[0\]\[5\] _2223_ _2209_ _2242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7157__A1 net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6879_ _2185_ _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8354__B1 _3527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8618_ _3173_ _3809_ _3810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8549_ _3716_ _3713_ _3714_ _3745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8657__A1 _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8409__A1 _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8682__B _3839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7396__A1 _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9088__CLK clknet_leaf_26_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7148__A1 _4362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6221__I _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8648__A1 _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6123__A2 _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7052__I _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7623__A2 _2868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8820__A1 _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5634__A1 _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7920_ _2736_ _3156_ _3158_ _3159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7851_ _3088_ _3091_ _3092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_110_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6802_ _2119_ _2088_ _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_64_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7782_ _2843_ _3024_ _3025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4994_ _4247_ _0436_ _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6733_ _2049_ _2052_ _2053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7139__A1 _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6664_ _1983_ _1984_ _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8403_ _3544_ _3603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5615_ _0890_ _0902_ _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6595_ _4263_ _1811_ _1917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5165__A3 _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8334_ _3517_ _3535_ _3536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5546_ _0981_ _0947_ _0929_ _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8265_ _3468_ _4272_ _3469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7311__A1 _2534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5477_ _0914_ _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7216_ _4095_ _2485_ _2484_ _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4428_ _4008_ _4009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_132_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7862__A2 _3102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8196_ _1602_ _3383_ _3415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_87_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4676__A2 _4098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5873__A1 _4073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7147_ _1444_ _2418_ _2419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8811__A1 _2307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7078_ _2342_ _2357_ _2358_ _1471_ _0165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6029_ _1217_ _1259_ _1262_ _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6050__A1 _4038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_3_0_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout52 net33 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4600__A2 _4159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8521__I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8948__CLK clknet_leaf_34_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7550__A1 _2298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5400__I1 as2650.r123_2\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8677__B _3856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6976__I _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7302__A1 _4090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7853__A2 _3087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4496__I _4076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7605__A2 _2851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8802__A1 _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5092__A2 _4021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8030__A2 _3263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5919__A2 _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_as2650_90 io_oeb[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XFILLER_127_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6592__A2 _1837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7475__C _2724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5400_ as2650.r123\[0\]\[7\] as2650.r123_2\[0\]\[7\] _4009_ _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6380_ as2650.stack\[3\]\[2\] _1715_ _1725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_75_wb_clk_i clknet_3_0_0_wb_clk_i clknet_leaf_75_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_127_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5331_ _0746_ _0770_ _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5790__I _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9103__CLK clknet_leaf_13_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8050_ _0902_ _3283_ _3284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5262_ _4281_ _0701_ _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7001_ _2280_ _1548_ _2284_ _2291_ _2292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_69_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5855__A1 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5193_ _0627_ _0633_ _4179_ _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_60_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5607__A1 as2650.r123\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8952_ _0113_ clknet_leaf_59_wb_clk_i as2650.stack\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7903_ _3139_ _3141_ _3142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8883_ _0044_ clknet_leaf_51_wb_clk_i as2650.stack\[1\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7834_ _2869_ _3066_ _3075_ _2735_ _3076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_58_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6032__A1 _4145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7666__B _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7765_ _2830_ _3007_ _3008_ _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5965__I _4037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4977_ as2650.r123\[2\]\[4\] as2650.r123_2\[2\]\[4\] _0339_ _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7780__A1 _3021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6716_ _0845_ _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7385__C _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7696_ _0603_ _0531_ _2941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_32_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6647_ _1820_ _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6578_ _1878_ _1900_ _1901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_121_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4897__A2 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8317_ _3500_ _3501_ _3518_ _3519_ _3520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5529_ _4308_ _0880_ _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8088__A2 _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8248_ _2258_ _2382_ _3451_ _2264_ _3452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_69_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8179_ _1640_ _3395_ _3396_ _3402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5205__I _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8516__I _3459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output31_I net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4821__A2 _4400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8012__A2 _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5377__A3 _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7523__A1 _2732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8251__A2 _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5065__A2 _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4900_ _0338_ _0341_ _0343_ _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__8003__A2 _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5880_ _1274_ _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_94_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4831_ _4360_ _4410_ _4281_ _4411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7550_ _2298_ _2545_ _2798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4762_ _4335_ _4341_ _4342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6501_ _1241_ _1394_ _1248_ _1804_ _1824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_140_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7481_ _1765_ _2686_ _2729_ _2730_ _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4693_ _4264_ _4272_ _4273_ _4274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_105_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7514__B2 as2650.stack\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6432_ _1741_ _1759_ _1760_ as2650.stack\[2\]\[7\] _1744_ _1764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_135_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6363_ _0967_ _1592_ _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_127_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8102_ _1422_ _3331_ _3332_ _3333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5314_ _0593_ _4318_ _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9082_ _0243_ clknet_leaf_25_wb_clk_i net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7817__A2 _3058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6294_ as2650.stack\[5\]\[7\] _1616_ _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_114_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8033_ _2547_ _3268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_103_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5245_ _0683_ _0684_ _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8490__A2 _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6096__A4 _4335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5176_ _0322_ _0616_ _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_60_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8242__A2 _3438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8793__A3 _2996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8935_ _0096_ clknet_3_1_0_wb_clk_i as2650.r123\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8866_ _0027_ clknet_leaf_48_wb_clk_i as2650.stack\[5\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6005__A1 _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_3_5_0_wb_clk_i clknet_0_wb_clk_i clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_73_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7817_ _2891_ _3058_ _3059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8797_ _3961_ _3965_ _3966_ _3659_ _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__9167__I net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7748_ _2546_ _2991_ _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_61_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7505__A1 _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7679_ _2689_ _2896_ _2893_ _2915_ _2924_ _2925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_123_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_67_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8233__A2 _3440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5047__A2 _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7744__A1 _2987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4730__A1 _4310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5030_ _0337_ _0332_ _4319_ _4416_ _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4684__I _4153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8224__A2 _3383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6981_ _4046_ _2270_ _2271_ _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_20_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6786__A2 _2102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5932_ _4159_ _1318_ _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8720_ _0387_ _2493_ _3892_ _3893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8651_ _3223_ _3831_ _3832_ _3834_ _3835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_61_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5863_ _0938_ _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__7735__A1 _4094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7602_ _2846_ _2848_ _2849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__4549__A1 _4128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4814_ _4064_ _4248_ _4394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8582_ _3500_ _3775_ _3519_ _3776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_37_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6002__A4 _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5794_ _1195_ _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7533_ _1353_ _1547_ _2781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4745_ _4163_ _4145_ _4325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_108_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7464_ _2710_ _2713_ _2714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4676_ _4024_ _4098_ _4257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8160__A1 _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6415_ _1590_ _1746_ _1753_ _0107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7395_ _1578_ _2647_ _2611_ _2648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xoutput18 net18 io_oeb[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_134_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput29 net53 io_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_6346_ as2650.r123\[3\]\[0\] _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4721__A1 _4290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9065_ _0226_ clknet_leaf_40_wb_clk_i as2650.stack\[6\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6277_ as2650.pc\[5\] _1643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8016_ _4005_ _1219_ _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5228_ _0335_ _0563_ _0367_ _0465_ _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__7671__B1 _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4594__I _4174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5159_ _0599_ _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5029__A2 _4319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8918_ _0079_ clknet_leaf_33_wb_clk_i as2650.stack\[5\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8849_ _0010_ clknet_leaf_67_wb_clk_i as2650.r123\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6314__I _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5201__A2 _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_123_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6701__A2 _1966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5268__A2 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6465__A1 as2650.stack\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4571__S0 _4018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7965__A1 _3195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8390__A1 _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8390__B2 _3590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7764__B _2927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6940__A2 _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7256__S _2501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4530_ _4014_ _4022_ _4111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8142__A1 _2623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4679__I _4088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4461_ _4041_ _4042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8693__A2 _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6200_ _0349_ _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7180_ _1271_ _4089_ _1552_ _4123_ _2451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_113_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6131_ _1232_ _1369_ _1483_ _1494_ _1516_ _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6456__A1 as2650.stack\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5259__A2 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6062_ _1418_ _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5013_ _0448_ _0449_ _4356_ _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6208__A1 _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7256__I0 _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7939__B _2894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6964_ _4092_ _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5431__A2 _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8703_ _0939_ _2324_ _3876_ _3877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_34_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5915_ _1203_ _1301_ _1306_ _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7971__A4 _3140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7708__A1 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6895_ _2026_ _2192_ _2198_ _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5982__A3 _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6134__I _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8634_ as2650.stack\[4\]\[9\] _3823_ _3824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5846_ _4040_ _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7184__A2 _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8381__A1 _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8565_ _1106_ _3484_ _3759_ _3760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5973__I _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5777_ _1110_ _1180_ _1184_ _0038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_5_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4728_ _4289_ _4308_ _4309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7516_ _2764_ _2765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8496_ _1491_ _0735_ _3693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7447_ _1297_ _2697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4659_ _4203_ _4240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6695__A1 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7378_ as2650.cycle\[4\] _2633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6329_ _1687_ _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9117_ _0278_ clknet_leaf_66_wb_clk_i as2650.psl\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8436__A2 _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9048_ _0209_ clknet_leaf_39_wb_clk_i as2650.pc\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6998__A2 _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6472__C _1773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5369__B _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8372__A1 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6922__A2 _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8124__A1 _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4499__I _4039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8675__A2 _3854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5489__A2 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5110__A1 _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6219__I _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4464__A3 _4044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7938__A1 _2885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_29_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_29_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_36_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4962__I _4142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8060__B1 _3280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6610__A1 _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8854__CLK clknet_leaf_68_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5700_ as2650.stack\[3\]\[11\] _1111_ _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_95_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6680_ _1938_ _1956_ _2001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5631_ _1059_ _1060_ _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5177__A1 _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5177__B2 _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6913__A2 _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8350_ _3549_ _3550_ _3551_ _3552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5562_ _0986_ _0996_ _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7301_ _2558_ _2439_ _2559_ _2560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4513_ as2650.addr_buff\[6\] _4094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8281_ _3458_ _3485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5493_ _4306_ _0882_ _0889_ _0925_ _0930_ _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_89_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7232_ _2493_ _2494_ _2499_ _1465_ _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_132_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4444_ as2650.ins_reg\[6\] _4025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7163_ net54 _2428_ _2434_ _2435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_144_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8418__A2 _3598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7513__I _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6429__A1 _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6114_ _0527_ _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7094_ _0288_ _2094_ _2368_ as2650.r123\[2\]\[4\] _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_100_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6045_ _1416_ _1420_ _1425_ _1431_ _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5101__A1 _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5652__A2 _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7929__A1 _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5968__I _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7996_ _1434_ _2400_ _3225_ _3230_ _3231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5404__A2 _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6947_ _2238_ _2239_ _2241_ _0151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8354__A1 _3534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7157__A2 _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6878_ _1542_ _1850_ _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__8354__B2 _3537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8617_ _3169_ _3773_ _3171_ _3809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5168__A1 _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5829_ _4073_ _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6904__A2 _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4915__A1 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8548_ _2831_ _3723_ _3743_ _3744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8106__A1 _3328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6117__B1 _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8479_ _3673_ _3676_ _3677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_118_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6668__A1 _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5340__A1 _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8409__A2 _3603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7093__A1 _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8877__CLK clknet_leaf_58_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6840__A1 _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5878__I _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7396__A2 _2411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8593__A1 _3144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7148__A2 _2416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8345__A1 _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4906__A1 _4143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8648__A2 _2571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7320__A2 _2575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5882__A2 _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5634__A2 _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5788__I _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7850_ _3089_ _3090_ _3091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8584__A1 _3126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6801_ _2078_ _2119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__9032__CLK clknet_leaf_23_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7781_ _3020_ _3023_ _3024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_17_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4993_ _0346_ _0435_ _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_63_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6732_ _2050_ _2051_ _2052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7139__A2 _2409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8336__A1 _4391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6663_ _1945_ _1954_ _1984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8113__B _3269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8402_ _2559_ _3602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5614_ _1043_ _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6594_ _4230_ _1908_ _1829_ _1915_ _1916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_34_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8333_ _2783_ _2786_ _3533_ _3535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5545_ _0334_ _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8639__A2 _3820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8264_ _4262_ _3468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5476_ _0913_ _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7311__A2 _2352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7215_ _2323_ _2485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5322__A1 as2650.r0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4427_ as2650.psl\[4\] _4008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_8195_ as2650.stack\[7\]\[0\] _3413_ _3414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6287__C _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5873__A2 _4077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7146_ _0527_ _1451_ _1216_ _2417_ _1253_ _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_119_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7075__A1 _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7077_ net23 _2357_ _2358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8811__A2 _2517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5625__A2 _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6822__A1 _4223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6028_ _1362_ _1392_ _1397_ _1414_ _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_100_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7979_ _1548_ _3212_ _3214_ _2335_ _3215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6050__A2 _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8327__A1 _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout53 net29 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_126_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6889__A1 _1923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5561__A1 _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7302__A2 _4056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5313__A1 _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7066__A1 _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_80 io_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_91 io_oeb[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XANTENNA__6041__A2 _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8318__A1 _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7328__I _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5330_ _0750_ _0755_ _0769_ _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5292__B _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5261_ _0700_ _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7063__I _2343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7000_ _1426_ _2290_ _2291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5855__A2 _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5192_ _0495_ _0502_ _0493_ _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_9_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_44_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_96_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5607__A2 _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8951_ _0112_ clknet_leaf_59_wb_clk_i as2650.stack\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7902_ _3140_ _3141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5311__I as2650.r0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8882_ _0043_ clknet_leaf_46_wb_clk_i as2650.stack\[2\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8557__A1 _3464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8557__B2 _2256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7833_ _2793_ _3070_ _3072_ _3074_ _3075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_110_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6032__A2 _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7764_ _1696_ _2878_ _2927_ _3008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_52_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4976_ _0418_ _4021_ _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6715_ _0418_ _1936_ _2035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7695_ _0538_ _0420_ _2940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6142__I _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6646_ _0349_ _1855_ _1967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7682__B _2927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5543__A1 _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6577_ _1883_ _1899_ _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_69_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8316_ _3473_ _3519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5528_ as2650.r123\[0\]\[2\] _0963_ _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8247_ _1064_ _2394_ _2330_ _1437_ _3451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_65_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5459_ _0896_ _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_57_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8178_ as2650.stack\[6\]\[4\] _3393_ _3401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9078__CLK clknet_leaf_51_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7129_ as2650.halted _1465_ _1543_ _2401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_59_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8796__A1 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8548__A1 _2831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7220__A1 _4189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8915__CLK clknet_leaf_35_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7771__A2 _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8720__A1 _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7523__A2 _2734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7592__B _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5891__I _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6936__B _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7039__A1 _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4896__I0 as2650.r123\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8251__A3 _2416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6227__I _1597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8539__A1 _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_opt_2_0_wb_clk_i clknet_3_5_0_wb_clk_i clknet_opt_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8003__A3 _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4970__I _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4830_ _4368_ _4409_ _4410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7762__A2 _2995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5287__B _4252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4761_ _4337_ _4340_ _4341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_60_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6500_ _1822_ _1823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7480_ _1294_ _2730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4692_ _4112_ _4061_ _4273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8711__A1 _3344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5525__A1 as2650.r123\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6431_ _1649_ _1758_ _1763_ _0113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6362_ _1589_ _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4879__A3 _4236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7278__A1 _2430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5313_ _0669_ _0752_ _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8101_ _1951_ _0873_ _3332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9081_ _0242_ clknet_leaf_24_wb_clk_i net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6293_ _1656_ _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8032_ _3244_ _3261_ _3266_ _3267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5244_ _0626_ _0630_ _0638_ _0647_ _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_114_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7293__A4 _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4500__A2 _4031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5175_ _0615_ _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7521__I _2460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8778__A1 _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6137__I _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8938__CLK clknet_leaf_42_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8934_ _0095_ clknet_opt_2_0_wb_clk_i as2650.r123\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4654__I3 as2650.r123_2\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8865_ _0026_ clknet_leaf_58_wb_clk_i as2650.stack\[5\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5976__I _4101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4880__I _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7816_ _3054_ _3057_ _3058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_101_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8796_ _0905_ _3961_ _3966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7753__A2 _2836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7747_ _2986_ _2943_ _2989_ _2991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_123_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4959_ _0395_ _0397_ _0401_ _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7678_ _2823_ _2923_ _2924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_138_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7505__A2 _2733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8702__A1 _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6629_ _0561_ _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8769__A1 _3940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5886__I _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7744__A2 _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5755__A1 _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4730__A2 _4192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7680__A1 _2881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7680__B2 _2688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4494__A1 _4064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6235__A2 _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7432__A1 _2671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6980_ _4119_ _4118_ _1246_ _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_93_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5931_ _1317_ _4337_ _0298_ _0386_ _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__5796__I _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8650_ _4195_ _2350_ _3234_ _3833_ _3834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5862_ _1256_ _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7735__A2 _2809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7601_ _2785_ _2786_ _2847_ _2848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_107_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4549__A2 _4129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4813_ _4392_ _4393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8581_ _3120_ _3774_ _3775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5793_ _1044_ _1194_ _1084_ _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_124_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7532_ _2779_ _2780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7944__C _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4744_ _4137_ _4324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7499__A1 as2650.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7463_ _2711_ _2712_ _2713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4675_ _4201_ _4255_ _4256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8121__B _4101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8160__A2 _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6414_ _1599_ _1749_ _1752_ as2650.stack\[2\]\[0\] _1745_ _1753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_128_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7394_ _2646_ _2647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xoutput19 net19 io_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__4721__A2 _4294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6345_ _1698_ _1676_ _1699_ _1700_ _0090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_103_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6276_ _0590_ _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_9064_ _0225_ clknet_leaf_39_wb_clk_i as2650.stack\[6\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5227_ _0666_ _0667_ _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_8015_ as2650.carry _3249_ _3250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7671__B2 as2650.stack\[5\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5158_ _0594_ _0596_ _0598_ _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_69_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7423__A1 _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5089_ as2650.r123\[2\]\[5\] as2650.r123_2\[2\]\[5\] _4012_ _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_44_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9116__CLK clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8917_ _0078_ clknet_leaf_33_wb_clk_i as2650.stack\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8848_ _0009_ clknet_3_1_0_wb_clk_i as2650.r123\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5737__A1 _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8779_ _3935_ _3949_ _3950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7426__I _2675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8257__I _2571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7161__I _2265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4571__S1 _4019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7265__I1 _2526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_62_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7717__A2 _2931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8390__A2 _2586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6940__A3 _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7336__I _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8142__A2 _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6240__I _4230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4460_ as2650.ins_reg\[4\] _4041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6130_ _1498_ _1505_ _1515_ _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_125_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_28_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6456__A2 _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6061_ _1434_ _1447_ _1448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5012_ _4276_ _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_39_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6208__A2 _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7256__I1 _2519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6843__C _2158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6963_ _1445_ _2253_ _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__8116__B _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8702_ _1445_ _2317_ _3874_ _3875_ _3876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5914_ as2650.stack\[0\]\[10\] _1304_ _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7169__B1 _2439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6894_ as2650.r123_2\[1\]\[3\] _2189_ _2197_ _2198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_59_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7708__A2 _2433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8633_ _3818_ _3823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5845_ _1074_ _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7184__A3 _2452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8381__A2 _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8630__I _3819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8564_ _3093_ _3758_ _3759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5776_ as2650.stack\[2\]\[9\] _1183_ _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7515_ as2650.stack\[3\]\[1\] _1296_ _1191_ as2650.stack\[0\]\[1\] as2650.stack\[1\]\[1\]
+ _1175_ _2764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
X_4727_ _4307_ _4308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8495_ _1393_ _3572_ _2482_ _3692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_120_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8133__A2 _3004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6144__A1 _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7446_ as2650.stack\[4\]\[0\] _1194_ _2695_ as2650.stack\[5\]\[0\] _0915_ _2696_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_4658_ _4238_ _4239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7892__A1 _2891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7377_ _2589_ _1058_ _2590_ _2632_ _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4589_ _4027_ _4070_ _4170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_9116_ _0277_ clknet_leaf_45_wb_clk_i as2650.overflow vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6328_ as2650.pc\[4\] _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_103_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9047_ _0208_ clknet_leaf_30_wb_clk_i as2650.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6259_ _0415_ _1627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_67_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5407__B1 _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5958__A1 _4142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8026__B _3260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4630__A1 _4210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7156__I _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8124__A2 _3263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6135__A1 _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7883__A1 _3089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4697__A1 _4265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7938__A2 _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8060__A1 _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6610__A2 _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4621__A1 _4192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_69_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_69_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_52_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5630_ _4046_ _4051_ _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6374__A1 _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5561_ _0461_ _0871_ _0963_ _0995_ _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8115__A2 _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7300_ _2409_ _2559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4512_ as2650.addr_buff\[7\] _4093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6126__A1 _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8280_ _3483_ _3484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5492_ _0929_ _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7874__A1 _3062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7231_ _2495_ _2496_ _2497_ _2498_ _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_4443_ _4023_ _4024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7162_ _2433_ _2434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6113_ net3 _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_113_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6429__A2 _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7093_ _0461_ _2361_ _2369_ _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6044_ _1426_ _1430_ _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7669__C _2470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7929__A2 _3141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8051__A1 _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7995_ _1093_ _1437_ _3227_ _3229_ _3230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_81_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6601__A2 _1922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6946_ _1000_ _2231_ _2214_ _2240_ _2241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_35_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6877_ _1698_ _2178_ _2184_ _0138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_70_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8616_ _3537_ _3804_ _3807_ _3763_ _2620_ _3808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_126_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5828_ _1222_ _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5168__A2 _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8547_ _3051_ _3558_ _3738_ _3742_ _3743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_124_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5759_ _1133_ _1164_ _1170_ _0034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4915__A2 _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6117__A1 _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8478_ _3634_ _3674_ _3675_ _3676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_118_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6117__B2 _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7865__A1 _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7429_ _1437_ _2331_ _2678_ _2679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_68_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7865__B2 _3105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5340__A2 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7617__A1 _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5224__I as2650.r0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7093__A2 _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4851__A1 as2650.holding_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8593__A2 _3766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6055__I _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4603__A1 _4162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8203__C _3409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4906__A2 _4099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8648__A3 _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6939__B _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7614__I _2860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5882__A3 _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8820__A3 _3911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4973__I as2650.r0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6831__A2 _2069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6800_ _2113_ _2117_ _2118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8971__CLK clknet_leaf_35_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7780_ _3021_ _3022_ _3023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6595__A1 _4263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4992_ _0433_ _0434_ _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6731_ _1942_ _1981_ _1998_ _2051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7139__A3 _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6662_ _1948_ _1953_ _1983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8401_ _2887_ _3600_ _3601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_31_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6898__A2 _2192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5613_ as2650.psu\[2\] _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6593_ _4379_ _1909_ _1914_ _1842_ _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_125_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8332_ _2783_ _3533_ _2786_ _3534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_30_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5544_ _0975_ _0979_ _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8263_ _1398_ _3466_ _3467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_118_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5475_ _0909_ _0912_ _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_132_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7311__A3 _2568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7214_ _1445_ _2480_ _2395_ _2483_ _2484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
X_4426_ _4006_ _4007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5322__A2 _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8194_ _3412_ _3413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_47_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7145_ _1074_ _1070_ _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_98_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5044__I _4325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8272__A1 _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7075__A2 _2355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7076_ _2347_ _2351_ _2352_ _2356_ _2357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_80_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5625__A3 _4119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6027_ _1396_ _1408_ _1413_ _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_104_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8575__A2 net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7978_ _2464_ _3213_ _1335_ _3214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5928__B _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6929_ _2220_ _2222_ _2226_ _0148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8327__A2 _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout54 net26 net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6889__A2 _2192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5010__A1 _4264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7838__A1 _3053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7838__B2 _2462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7434__I _2683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8844__CLK clknet_leaf_69_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6510__A1 _4279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8263__A1 _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7066__A2 _2344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5077__A1 _4012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5889__I _4109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4824__A1 _4252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8015__A1 as2650.carry vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_70 io_oeb[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7774__B1 _2956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_as2650_81 io_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xwrapped_as2650_92 io_oeb[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_2673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5001__A1 _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5552__A2 _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5292__C _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5260_ _0622_ _0682_ _0697_ _0699_ _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XANTENNA__6501__A1 _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5191_ _0385_ _0631_ _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8254__A1 _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5799__I _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8950_ _0111_ clknet_leaf_34_wb_clk_i as2650.stack\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7901_ _3111_ _3084_ _3140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8006__A1 _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8881_ _0042_ clknet_leaf_47_wb_clk_i as2650.stack\[2\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_13_wb_clk_i clknet_3_2_0_wb_clk_i clknet_leaf_13_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_92_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7832_ _1578_ _3058_ _3073_ _1248_ _3074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_64_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6568__A1 _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6032__A3 _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7763_ _2968_ _2977_ _3006_ _2688_ _3007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4975_ _0417_ _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6714_ _2032_ _2033_ _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7694_ _1644_ _2938_ _2939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_36_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6645_ _1917_ _1966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6576_ _1885_ _1898_ _1899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__8867__CLK clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6740__A1 _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8315_ _3463_ _3494_ _3516_ _3517_ _3518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_117_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_3_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5527_ _0877_ _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8246_ _2419_ _2423_ _3449_ _3450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_69_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5458_ as2650.psu\[1\] _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_121_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8177_ _1727_ _3398_ _3399_ _3400_ _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_99_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5389_ _0826_ _0827_ _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8245__A1 _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7128_ _4301_ _4084_ _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5059__A1 _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7203__B _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7059_ _4166_ _2337_ _2340_ _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5502__I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6559__A1 _4209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7220__A2 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output17_I net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5231__A1 _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5782__A2 _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8720__A2 _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6731__A1 _1942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5534__A2 _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4788__I _4367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9022__CLK clknet_leaf_7_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7039__A2 _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8787__A2 _3951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6444__S _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6243__I _1612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4760_ _4175_ _4338_ _4339_ _4340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5773__A2 _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7783__B _2489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4691_ _4271_ _4272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6430_ _1651_ _1759_ _1760_ as2650.stack\[2\]\[6\] _1744_ _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__5525__A2 _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6361_ _1708_ _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8100_ _3253_ _2923_ _3330_ _0935_ _3331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5312_ _0751_ _4415_ _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8475__A1 _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7278__A2 _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9080_ _0241_ clknet_leaf_65_wb_clk_i as2650.stack\[7\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6292_ _1655_ _1656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8031_ _1580_ _4250_ _3265_ _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5243_ as2650.holding_reg\[6\] _0599_ _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_88_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5174_ _0582_ _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8119__B _3348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8778__A2 _3920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6418__I _1744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7958__B _2948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8933_ _0094_ clknet_leaf_75_wb_clk_i as2650.r123\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8864_ _0025_ clknet_leaf_53_wb_clk_i as2650.stack\[5\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_36_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7815_ _2974_ _3055_ _3056_ _3057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6005__A3 _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8795_ _2832_ _3962_ _3964_ _3920_ _3965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_52_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7746_ _2986_ _2943_ _2989_ _2990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4958_ _4129_ _0400_ _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7677_ _0923_ _2916_ _2917_ _2922_ _2923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_138_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4889_ _0332_ _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_71_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8702__A2 _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6628_ _1946_ _1949_ _1950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_137_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6713__A1 _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9045__CLK clknet_leaf_29_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6559_ _4209_ _4416_ _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9116__D _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8229_ _1190_ _3437_ _3439_ _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8218__A1 _1738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8769__A2 _3938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7977__B1 _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7868__B _2927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7159__I _2430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4638__S0 _4003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6063__I _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5755__A2 _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6704__A1 _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9026__D _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8457__A1 _2791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7665__C1 _2890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8209__A1 _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4494__A2 _4074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6235__A3 _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5930_ _4293_ _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_47_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5861_ _1255_ _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7196__A1 _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7600_ _1621_ _1402_ _2847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4812_ _4391_ _4392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8580_ _3123_ _3773_ _3774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6943__A1 as2650.r123_2\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5792_ _1193_ _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7531_ _2778_ _2779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__9068__CLK clknet_leaf_42_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4743_ _4138_ _4283_ _4305_ _4323_ _0000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_109_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7499__A2 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8696__A1 _3869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7462_ _1596_ _4242_ _2712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4674_ _4205_ _4224_ _4254_ _4255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6413_ _1751_ _1752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7393_ _2430_ _1334_ _2646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_128_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6344_ _1657_ _1680_ _1681_ _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_1_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4721__A3 _4301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_9063_ _0224_ clknet_leaf_37_wb_clk_i as2650.stack\[6\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7120__A1 _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8905__CLK clknet_leaf_62_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6275_ _1636_ _1637_ _1641_ _0079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7532__I _2779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8014_ _3248_ _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5226_ _0564_ _0665_ _0561_ _0525_ _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__7671__A2 _2692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5157_ _4218_ _0597_ _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7423__A2 _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8620__A1 _2898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5088_ _0519_ _0522_ _0526_ _0529_ _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5987__I _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5434__A1 _4004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4891__I as2650.r0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8916_ _0077_ clknet_leaf_33_wb_clk_i as2650.stack\[5\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7187__A1 _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8847_ _0008_ clknet_leaf_67_wb_clk_i as2650.r123\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5737__A2 _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8778_ _1572_ _3920_ _3949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_90_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7729_ _1643_ _0603_ _2972_ _2973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5936__B _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8687__A1 _3851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8439__A1 _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7111__A1 _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7442__I _2691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8611__A1 _3595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7414__A2 _2355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5425__A1 _4111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6925__A1 _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7350__A1 _2550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8928__CLK clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5581__B _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7102__A1 _4005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6060_ _1435_ _1437_ _1441_ _1446_ _1447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input8_I io_in[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5011_ _4277_ _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8602__A1 _3147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6208__A3 _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7301__B _2559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7956__A3 _3141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6962_ _1846_ _1543_ _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_4_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5913_ _1200_ _1301_ _1305_ _0053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8701_ _1464_ _1544_ _3875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7169__A1 _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6893_ _0483_ _2012_ _2197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7169__B2 net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8632_ _1190_ _3820_ _3822_ _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_62_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5844_ _1230_ _1238_ _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6916__A1 _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8563_ _1106_ _3525_ _3757_ _3654_ _2437_ _3758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_107_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5775_ _1178_ _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7527__I _2684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7514_ as2650.stack\[7\]\[1\] _2762_ _1046_ as2650.stack\[6\]\[1\] _0913_ _2763_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__8669__A1 _3836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4726_ _4291_ _4307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8494_ _3688_ _3689_ _3690_ _3691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_120_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7445_ _2694_ _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7341__A1 _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6144__A2 _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4657_ _4237_ _4238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7376_ _2591_ _2619_ _2631_ _2589_ _2632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__7892__A2 _3125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4588_ _4157_ _4169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9115_ _0276_ clknet_leaf_42_wb_clk_i as2650.psu\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6327_ _1629_ _1662_ _1686_ _0086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9046_ _0207_ clknet_leaf_40_wb_clk_i as2650.pc\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_67_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6258_ _1620_ _1595_ _1626_ _0077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_130_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5209_ _0649_ _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6189_ _1559_ _1565_ _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8093__I _2594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5510__I _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5958__A2 _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6080__A1 _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7437__I _2437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6135__A2 _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5894__A1 _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8268__I _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4796__I _4375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7096__B1 _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8832__A1 _2518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4449__A2 as2650.cycle\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5646__A1 _4003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6446__I0 _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8060__A2 _3276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6071__A1 _4109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4621__A2 _4077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6374__A2 _1712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6251__I _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5560_ _0415_ _0882_ _0889_ _0994_ _0930_ _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_106_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_38_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4511_ _4091_ _4092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7791__B _3033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5491_ _4309_ _0928_ _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6126__A2 _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7230_ _4194_ _1454_ _2498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9106__CLK clknet_leaf_13_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4442_ _4017_ _4022_ _4023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7874__A2 _3097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4688__A2 as2650.addr_buff\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5885__A1 _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_37_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7161_ _2265_ _2433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7087__B1 _2364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6112_ _1484_ _1495_ _0536_ _0605_ _1497_ _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__7626__A2 _2871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8823__A1 _3978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7092_ _0288_ _2054_ _2368_ as2650.r123\[2\]\[3\] _2369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5637__A1 _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6043_ _1429_ _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7994_ _4133_ _2676_ _2276_ _3228_ _3229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_113_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6945_ _1008_ _2218_ _2240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6876_ _1741_ _2179_ _2180_ as2650.stack\[0\]\[7\] _2165_ _2184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_8615_ net40 _3806_ _3807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_50_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5827_ _1073_ _4099_ _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_76_wb_clk_i_I clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8546_ _3740_ _3741_ _2458_ _3742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5758_ as2650.stack\[6\]\[12\] _1166_ _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4709_ _4289_ _4290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8477_ _3639_ _0618_ _3675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_108_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6117__A2 _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5689_ as2650.r123\[0\]\[2\] _1113_ _1116_ _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_68_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7428_ _2676_ _2677_ _1561_ _2678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__7865__A2 _2961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7206__B _1563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4923__I0 as2650.r123\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7359_ _2613_ _2614_ _2615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_85_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7617__A2 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9029_ _0190_ clknet_leaf_17_wb_clk_i as2650.cycle\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4851__A2 _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5240__I _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4603__A2 _4165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7167__I _4194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8500__B _3464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7305__A1 _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9034__D _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7608__A2 _2853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8805__A1 _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8805__B2 _3973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5619__A1 _4141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6246__I _1606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5150__I _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6044__A1 _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4991_ _0304_ _4398_ _0294_ _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__7792__A1 _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6595__A2 _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6730_ _1985_ _1997_ _2050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6661_ _1942_ _1981_ _1982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8400_ _2844_ _3599_ _3600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5612_ _1038_ _1042_ _0015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5555__B1 _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6592_ _0355_ _1837_ _1838_ _1913_ _1914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_8331_ as2650.pc\[0\] net5 _2748_ _3533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5543_ _0916_ _0976_ _0978_ _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_129_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8262_ _3465_ _4279_ _3466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7847__A2 _2987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5474_ _0910_ _0911_ _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7213_ _2481_ _1552_ _2482_ _2325_ _2483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_105_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7311__A4 _2569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4425_ _4005_ _4006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8193_ _3411_ _3412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7144_ _2415_ _2416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4530__A1 _4014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8272__A2 _2897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7075_ _2354_ _2355_ _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6026_ _1411_ _1287_ _1412_ _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_101_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5625__A4 _4033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7783__A1 _2599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7977_ _4094_ _2861_ _2445_ _3208_ _2433_ _3213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6928_ as2650.r123_2\[0\]\[1\] _2224_ _2225_ _2210_ _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_126_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7535__A1 as2650.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6859_ _1670_ _2169_ _2171_ as2650.stack\[0\]\[1\] _2166_ _2173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_17_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5010__A2 _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8529_ _3667_ _3669_ _3724_ _3687_ _3725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_136_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5849__A1 _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5077__A2 as2650.r123\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6274__A1 _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6274__B2 as2650.stack\[5\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4824__A2 _4390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8015__A2 _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6026__A1 _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xwrapped_as2650_60 io_oeb[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_3386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7774__A1 as2650.stack\[4\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_as2650_71 io_oeb[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__8281__I _3458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7774__B2 as2650.stack\[5\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_as2650_82 io_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_93 io_oeb[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7526__A1 _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4760__A1 _4175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6501__A2 _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5190_ _0627_ _0630_ _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_79_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4984__I _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6265__A1 as2650.stack\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4917__C _4198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4815__A2 _4249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7900_ as2650.pc\[11\] _3139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_95_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8880_ _0041_ clknet_leaf_47_wb_clk_i as2650.stack\[2\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7831_ _1577_ _3053_ _3073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4933__B _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7765__A1 _2830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8191__I _3409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7762_ _2976_ _2995_ _3005_ _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4974_ _0416_ _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_53_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_53_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_71_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6713_ _1989_ _1996_ _2033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7693_ _1638_ _2907_ _2938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7517__A1 as2650.stack\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6644_ _1856_ _1965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6575_ _1890_ _1897_ _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_121_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8314_ _2409_ _3517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5526_ _0945_ _4136_ _4412_ _0962_ _0009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__4751__A1 _4178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8245_ _2402_ _3448_ _3449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5457_ _0894_ _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4503__A1 _4080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8176_ _1729_ _3395_ _3396_ _3400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5388_ _0710_ _4321_ _0753_ _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_120_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7127_ _1554_ _1546_ _2397_ _2398_ _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_141_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5059__A2 _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7058_ net22 _2337_ _2339_ _2340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6009_ _1395_ _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8315__B _3516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6559__A2 _4416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7756__A1 _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6614__I _1935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5231__A2 _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7508__A1 _2744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8705__B1 _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5519__B1 _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4990__A1 _4076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4742__A1 _4306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8961__CLK clknet_leaf_56_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8276__I _3479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8236__A2 _3437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7995__A1 _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6460__S _1778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4981__A1 _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4690_ _4265_ _4270_ _4271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__8172__A1 _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6722__A2 _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6360_ as2650.r123\[3\]\[7\] _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5311_ as2650.r0\[5\] _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8475__A2 _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6291_ as2650.pc\[7\] _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_66_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6486__A1 _4098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5289__A2 _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8030_ _3262_ _3263_ _3264_ _1559_ _3265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_88_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5242_ as2650.holding_reg\[6\] _0681_ _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_130_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5173_ _4368_ _0613_ _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6238__A1 _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8119__C _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6238__B2 as2650.stack\[5\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7986__A1 _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6789__A2 _2106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput1 io_in[10] net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8932_ _0093_ clknet_leaf_73_wb_clk_i as2650.r123\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7958__C _3039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8863_ _0024_ clknet_leaf_54_wb_clk_i as2650.stack\[5\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7738__A1 _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7738__B2 _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6434__I _1667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7814_ _1794_ _1737_ _0724_ _3056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_91_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8794_ _0905_ _3963_ _3964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7745_ _2988_ _2989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_40_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4957_ _0399_ _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_36_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8789__C _3659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4888_ _4382_ _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7676_ as2650.stack\[2\]\[4\] _2692_ _2919_ _2921_ _2922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_138_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8702__A3 _3874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6627_ _0416_ _0524_ _1949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8984__CLK clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4724__A1 as2650.r123\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6558_ _0838_ _1879_ _1880_ _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_106_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5509_ _0941_ _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6489_ _4082_ _1811_ _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6477__A1 _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7674__B1 _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8228_ as2650.stack\[7\]\[8\] _3438_ _3439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8218__A2 _3412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8159_ _3385_ _3386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5513__I _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7977__A1 _4094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7977__B2 _3208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7029__I0 _2312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4638__S1 _4014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6952__A2 _2243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8154__A1 _3372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4799__I _4249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7175__I _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4715__A1 _4131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8457__A2 _2936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7665__B1 _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7665__C2 _2710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6519__I _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5140__A1 _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5423__I _4110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5691__A2 _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7968__A1 _2591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8090__B1 _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6640__A1 _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8857__CLK clknet_leaf_57_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6254__I _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5860_ _1254_ _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8393__A1 net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4811_ net6 _4391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5791_ _1192_ _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7530_ _2539_ _2706_ _2778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4742_ _4306_ _4317_ _4322_ _4323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_109_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8145__A1 _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7461_ as2650.pc\[0\] net5 _2711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4673_ _4228_ _4239_ _4240_ _4253_ _4254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__8696__A2 _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6412_ _1713_ _0973_ _1750_ _1751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4502__I _4082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7392_ _2641_ _2642_ _2644_ _2645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_122_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6343_ as2650.stack\[4\]\[7\] _1677_ _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6459__A1 _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9062_ _0223_ clknet_leaf_38_wb_clk_i as2650.stack\[6\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6274_ _1640_ _1625_ _1607_ as2650.stack\[5\]\[4\] _1608_ _1641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_131_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7120__A2 _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5225_ _0564_ _0561_ _0525_ _0665_ _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8013_ _3247_ _3248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_9_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5156_ as2650.r123\[1\]\[6\] as2650.r123\[0\]\[6\] as2650.r123_2\[1\]\[6\] as2650.r123_2\[0\]\[6\]
+ _4003_ _4013_ _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_57_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7969__B _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8620__A2 _3807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5087_ _0527_ _0528_ _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_84_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5434__A2 _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8915_ _0076_ clknet_leaf_35_wb_clk_i as2650.stack\[5\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7974__A4 _3155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8846_ _0007_ clknet_leaf_69_wb_clk_i as2650.r123\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7187__A2 _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8384__A1 _2788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_77_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8777_ _3936_ _3947_ _3948_ _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_40_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5989_ _1375_ _1374_ _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7728_ _2933_ _2971_ _2972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4945__A1 _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8136__A1 _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8687__A2 _3863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7659_ _1410_ _2593_ _2905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5508__I _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6698__A1 _2014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7647__B1 _2890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7111__A2 _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6339__I _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6870__A1 _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8072__B1 _3302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6622__A1 _1942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5425__A2 _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7178__A2 _4122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8375__A1 _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_44_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6925__A2 _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8127__A1 _3338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8222__C _3408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8678__A2 _3846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7350__A2 _2606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_4_0_wb_clk_i clknet_0_wb_clk_i clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_67_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7102__A2 _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5113__A1 _4367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5010_ _4264_ _0452_ _4273_ _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_79_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6961_ as2650.addr_buff\[0\] _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_47_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9035__CLK clknet_leaf_40_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8700_ _0403_ _1846_ _3874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5912_ as2650.stack\[0\]\[9\] _1304_ _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_81_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7169__A2 _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8366__A1 _3540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6892_ _1979_ _2186_ _2195_ _2196_ _0141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_59_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8631_ as2650.stack\[4\]\[8\] _3821_ _3822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5843_ _1231_ _1237_ _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8562_ _2862_ _3754_ _3098_ _3757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_66_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5774_ _1103_ _1180_ _1182_ _0037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8132__C _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7513_ _0911_ _2762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8669__A2 _3849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4725_ _4189_ _4306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8493_ _3688_ _3689_ _3572_ _3690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7444_ _1175_ _2694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4656_ _4232_ _4234_ _4236_ _4237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__7341__A2 _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6144__A3 _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7375_ _2621_ _2628_ _2630_ _2326_ _2631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_116_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7543__I _2460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4587_ _4167_ _4168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9114_ _0275_ clknet_leaf_44_wb_clk_i as2650.psu\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6326_ as2650.stack\[4\]\[3\] _1665_ _1685_ _1660_ _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_107_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5104__A1 _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9045_ _0206_ clknet_leaf_29_wb_clk_i as2650.pc\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6257_ _1624_ _1625_ _1607_ as2650.stack\[5\]\[2\] _1608_ _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_89_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5655__A2 _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5208_ _0622_ _0625_ _0645_ _0648_ _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_88_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6188_ _1564_ _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5998__I _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_131_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5139_ _0323_ _0300_ _0398_ _0424_ _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_96_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6604__A1 _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5958__A3 _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_8_wb_clk_i clknet_3_2_0_wb_clk_i clknet_leaf_8_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_26_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6080__A2 _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8357__A1 _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8829_ _2525_ _3992_ _1492_ _3994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6907__A2 _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4918__A1 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8109__A1 _3324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6135__A3 _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5343__A1 _4206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5894__A2 _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7096__A1 _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8293__B1 _3493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6843__A1 _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5646__A2 _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9058__CLK clknet_leaf_39_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8596__A1 _3143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6446__I1 as2650.stack\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6071__A2 _4225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8348__A1 _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4909__A1 _4039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5148__I _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4510_ _4090_ _4055_ _4091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5490_ _0879_ _0927_ _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7323__A2 _2564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4987__I _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4441_ _4021_ _4022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_78_wb_clk_i clknet_3_0_0_wb_clk_i clknet_leaf_78_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5885__A2 _4308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7160_ _4070_ _1348_ _1460_ _2431_ _2432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_67_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7087__A1 _4317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6111_ _1496_ _4249_ _1497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7091_ _2363_ _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6042_ _1428_ _4125_ _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5637__A2 _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8194__I _3412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8587__A1 _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6598__B1 _1916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7993_ _2652_ _2673_ _3228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_81_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6944_ _2067_ _2229_ _2239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8143__B _3324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6875_ _1649_ _2178_ _2183_ _0137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_74_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8614_ _3805_ _3791_ _3806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5486__C _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5826_ _1215_ _1220_ _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_23_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8545_ _3054_ _3739_ _2629_ _3741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5573__A1 _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5757_ _1126_ _1163_ _1169_ _0033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8797__C _3659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4708_ _4286_ _4288_ _4289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_135_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8476_ _3639_ _0618_ _3674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__8511__A1 _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5688_ _1115_ _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_108_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7427_ _1450_ _1091_ _2677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4639_ _4218_ _4219_ _4220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7358_ _1054_ _1247_ _1058_ _2614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7206__C _2476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4923__I1 as2650.r123_2\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5007__B _4371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6309_ _0967_ _1602_ _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8814__A2 _3911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7289_ _4081_ _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_77_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6825__A1 _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9028_ _0189_ clknet_leaf_17_wb_clk_i as2650.cycle\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8578__A1 _3763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7250__A1 _1627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8918__CLK clknet_leaf_33_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8053__B _4078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7002__A1 _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7553__A2 _2799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8502__A1 net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5316__A1 _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5867__A2 _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7069__A1 _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8805__A2 _3969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5619__A2 _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9050__D _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8569__A1 _3472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6971__B _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6044__A2 _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7241__A1 _4326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6463__S _1778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4990_ _4076_ _0323_ _0301_ _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__7792__A2 _2991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6660_ _1941_ _1944_ _1981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7544__A2 _2790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8741__A1 _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5611_ _0817_ _0869_ _0946_ _1041_ _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5555__A1 as2650.stack\[2\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5555__B2 as2650.stack\[0\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6591_ _1400_ _1910_ _1912_ _1821_ _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_8330_ _3531_ _3532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5542_ as2650.stack\[7\]\[10\] _0977_ _0969_ as2650.stack\[6\]\[10\] _0978_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_9_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7307__B _2560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5307__A1 _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8261_ _4365_ _3465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5473_ _0894_ _0896_ _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7212_ _2255_ _2482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4424_ _4004_ _4005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8192_ _1146_ _0900_ _1605_ _3411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_144_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7143_ _1056_ _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7821__I _3062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6807__A1 _2071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7074_ _1069_ _2318_ _2355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_140_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6025_ _1374_ _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_45_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7232__A1 _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8652__I _3835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7976_ _3038_ _2979_ _3211_ _3029_ _3212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7783__A2 _3011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6927_ _1922_ _2208_ _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6172__I _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6858_ _1590_ _2167_ _2172_ _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7535__A2 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8732__A1 _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5809_ _1132_ _1207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5546__A1 _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6789_ _1964_ _2106_ _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8528_ _0783_ _0780_ _3724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8459_ net33 _3488_ _3658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5516__I _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5849__A2 _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4420__I as2650.ins_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8827__I _3991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8799__A1 _1859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7887__B _3126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7223__A1 _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6026__A2 _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_61 io_oeb[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_as2650_72 io_oeb[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_3398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8890__CLK clknet_leaf_41_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_as2650_83 io_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5785__A1 _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_94 io_oeb[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_2686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7526__A2 _2731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8723__A1 _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5001__A3 _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6501__A3 _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5161__I _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7214__A1 _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7830_ _3063_ _2861_ _3071_ _1398_ _1353_ _3072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__8411__B1 _3549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7761_ _2996_ _2968_ _3004_ _2823_ _3005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__5776__A1 as2650.stack\[2\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4973_ as2650.r0\[4\] _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6712_ _1991_ _1995_ _2032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7692_ _2782_ _2931_ _2936_ _2603_ _2937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7517__A2 _2691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8714__A1 _3869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5528__A1 as2650.r123\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6643_ _1963_ _1964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6574_ _1893_ _1896_ _1897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8313_ _3508_ _3514_ _3515_ _3516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5525_ as2650.r123\[0\]\[1\] _0942_ _0961_ _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4751__A2 _4167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8244_ _2675_ _1561_ _2665_ _1050_ _3448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5456_ as2650.psu\[0\] _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_86_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8175_ as2650.stack\[6\]\[3\] _3393_ _3399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5387_ _0588_ _4417_ _0670_ _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_114_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7126_ _4108_ _1219_ _2398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6167__I _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7057_ _2338_ _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__9119__CLK clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6008_ _1394_ _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7205__A1 _2462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_110_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7959_ _1129_ _1121_ _3155_ _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8705__A1 _4207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8705__B2 _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4990__A2 _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8181__A2 _3393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4742__A2 _4317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7692__A1 _2782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6077__I _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7995__A2 _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7636__I _2707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5310_ _0663_ _0673_ _0749_ _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6290_ _1653_ _1654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7683__A1 _2830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6486__A2 _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5241_ _0680_ _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4497__A1 _4073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5172_ _4370_ _0587_ _0612_ _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_111_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7986__A2 _4081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput2 io_in[11] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_133_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8931_ _0092_ clknet_3_4_0_wb_clk_i as2650.r123\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5997__A1 _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8416__B _3515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8862_ _0023_ clknet_leaf_49_wb_clk_i as2650.stack\[5\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7738__A2 _2968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7813_ _2969_ _3020_ _3055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_37_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8793_ _0881_ _3940_ _2996_ _3963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_52_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7744_ _2987_ _0595_ _2988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_40_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4956_ _0398_ _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7675_ _2920_ _2921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_123_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4887_ _0330_ _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6626_ _0849_ _1946_ _1947_ _1894_ _1948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_14_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5921__A1 _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4724__A2 _4304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6557_ _0837_ _0840_ _1880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_14_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5508_ _0860_ _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6488_ _4310_ _1095_ _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8227_ _3436_ _3438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6477__A2 _4314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5439_ _4017_ _0876_ _0870_ _4285_ _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7674__B2 as2650.stack\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8158_ _3384_ _3385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6229__A2 _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7109_ _1341_ _4170_ _1235_ _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_82_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8089_ _1580_ _0436_ _3320_ _3321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7977__A2 _2861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9091__CLK clknet_leaf_25_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7029__I1 _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7729__A2 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8045__C _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output22_I net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4715__A2 _4295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_17_wb_clk_i_I clknet_opt_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8287__I _3483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7665__A1 as2650.addr_buff\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7665__B2 _2881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5140__A2 _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7417__A1 _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8090__A1 _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5979__A1 _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6640__A2 _1923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4651__A1 _4230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4810_ _4389_ _4390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5790_ _1191_ _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_56_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4741_ _4321_ _4322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7366__I _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7460_ _1240_ _1443_ _2710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4672_ _4243_ _4246_ _4251_ _4252_ _4253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_135_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6411_ _1082_ _1750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7391_ _1843_ _2643_ _2611_ _2644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6342_ _1653_ _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_127_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6459__A2 _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9061_ _0222_ clknet_leaf_38_wb_clk_i as2650.stack\[6\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6273_ _1639_ _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_103_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7120__A3 _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8012_ _4004_ _1218_ _3247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5224_ as2650.r0\[0\] _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7408__A1 _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5155_ _4214_ _0595_ _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5086_ _4019_ _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8914_ _0075_ clknet_leaf_33_wb_clk_i as2650.stack\[5\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8845_ _0006_ clknet_leaf_69_wb_clk_i as2650.r123\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8384__A2 _2849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8951__CLK clknet_leaf_59_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8776_ _1747_ _3936_ _2534_ _3948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6395__A1 _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5988_ as2650.psl\[6\] _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7727_ as2650.pc\[5\] net1 _2971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4939_ as2650.holding_reg\[3\] _0344_ _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4945__A2 _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8136__A2 _4223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6147__A1 _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7209__C _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7658_ _2900_ _2865_ _2902_ _2904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_123_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7895__A1 _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6609_ _1881_ _1882_ _1931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__7895__B2 _2832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7589_ _2819_ _2836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_opt_1_0_wb_clk_i clknet_3_3_0_wb_clk_i clknet_opt_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_21_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7647__A1 _2885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7647__B2 _2892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4881__A1 _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8072__A1 _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8375__A2 _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6386__A1 _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6138__A1 _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5361__A2 _4222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9053__D _0214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7102__A3 _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5113__A2 _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8063__A1 _2623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8974__CLK clknet_leaf_57_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6960_ _1653_ _2231_ _2210_ _2251_ _0154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_81_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5911_ _1299_ _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6891_ _0380_ _2071_ _2196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8630_ _3819_ _3821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5842_ _0938_ _1236_ _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_107_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8561_ _3602_ _3747_ _3755_ _2459_ _3756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_37_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4927__A2 _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5773_ as2650.stack\[2\]\[8\] _1181_ _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5609__I _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7512_ as2650.stack\[4\]\[1\] _1193_ _2694_ as2650.stack\[5\]\[1\] _2761_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4724_ as2650.r123\[1\]\[0\] _4304_ _4305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6129__A1 _4005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8492_ _1519_ _0781_ _3689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7443_ as2650.stack\[7\]\[0\] _1298_ _2692_ as2650.stack\[6\]\[0\] _2693_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4655_ _4217_ _4235_ _4236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XFILLER_116_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7374_ _1523_ _2629_ _2410_ _2440_ _2630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5352__A2 _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4586_ _4166_ _4143_ _4167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7045__B _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7629__A1 _2834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9113_ _0274_ clknet_leaf_43_wb_clk_i as2650.psu\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6325_ _1684_ _1672_ _1685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5344__I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9044_ _0205_ clknet_leaf_29_wb_clk_i as2650.pc\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5104__A2 _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6256_ _1603_ _1625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8655__I _3835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5207_ _0299_ _0647_ _0622_ _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_131_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6187_ _1551_ _1563_ _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_57_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8054__A1 _3282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5138_ _4324_ _0558_ _0579_ _0004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6604__A2 _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5069_ _0510_ _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4615__A1 _4193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5958__A4 _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6080__A3 _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8357__A2 _3558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8828_ _1584_ _3952_ _2524_ _3993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_73_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8759_ _1273_ _1068_ _2467_ _3930_ _3931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_40_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8109__A2 _2096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4423__I _4003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5591__A2 _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7868__A1 _2685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6135__A4 _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8847__CLK clknet_leaf_67_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6540__A1 _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5343__A2 _4379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8293__A1 _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7096__A2 _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8293__B2 _3495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6843__A2 _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8045__A1 _3277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8596__A2 _2482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8348__A2 _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4909__A2 _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5582__A2 _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7859__A1 _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4440_ _4020_ _4021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5164__I _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6110_ net5 _1496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_98_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8284__A1 _3338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7087__A2 _1960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7090_ _0366_ _2361_ _2367_ _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9002__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6041_ _1427_ _1247_ _1428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4845__A1 _4324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_47_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_47_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_67_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8587__A2 _3480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4508__I _4088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7992_ _4363_ _3226_ _4260_ _2656_ _3227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__6598__A1 _4359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6943_ as2650.r123_2\[0\]\[4\] _2224_ _2227_ _2238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_78_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6874_ _1651_ _2179_ _2180_ as2650.stack\[0\]\[6\] _2165_ _2183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_81_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8613_ net39 _3805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_50_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5825_ _4006_ _1217_ _1219_ _1092_ _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_22_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8544_ _3054_ _3739_ _3740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5756_ as2650.stack\[6\]\[11\] _1166_ _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_72_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4707_ _4287_ _4284_ _4288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8475_ _0725_ _0734_ _3673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_33_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5687_ _1114_ _1089_ _1097_ as2650.r123_2\[0\]\[2\] _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_120_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8511__A2 _2862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7426_ _2675_ _2676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_120_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4638_ as2650.r123\[1\]\[7\] as2650.r123\[0\]\[7\] as2650.r123_2\[1\]\[7\] as2650.r123_2\[0\]\[7\]
+ _4003_ _4014_ _4219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_89_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7357_ _4029_ _4121_ _4103_ _2613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_78_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4569_ as2650.r123\[1\]\[0\] as2650.r123_2\[1\]\[0\] _4010_ _4150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7078__A2 _2357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8275__A1 _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6308_ _1614_ _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7288_ _2546_ _2547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9027_ _0188_ clknet_leaf_17_wb_clk_i as2650.cycle\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6825__A2 _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6239_ _1590_ _1595_ _1609_ _0075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_131_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6589__A1 _4106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5013__A1 _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8750__A2 _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8502__A2 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5316__A2 _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7710__B1 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9025__CLK clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8266__A1 _1496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7069__A2 _2349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8509__B _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8295__I _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5619__A3 _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8569__A2 _2286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8244__B _2665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4772__B _4164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7792__A3 _3033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5159__I _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5610_ _1040_ _4309_ _0882_ _0928_ _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__8741__A2 _3262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5555__A2 _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6590_ _4400_ _1911_ _1912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5541_ _0892_ _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8260_ _2287_ _3464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5307__A2 _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5472_ as2650.psu\[2\] _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6504__A1 _4239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7211_ _2267_ _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4423_ _4003_ _4004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8191_ _3409_ _3410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7142_ _0965_ _2406_ _2413_ _2414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_119_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7323__B _2580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6807__A2 _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7073_ _2353_ _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4818__A1 _4265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6024_ _1410_ _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5491__A1 _4309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7977__C _2433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7232__A2 _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7975_ as2650.pc\[14\] _3210_ _3211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8154__B _3276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6926_ _2223_ _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6857_ _1598_ _2169_ _2171_ as2650.stack\[0\]\[0\] _2166_ _2172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__5069__I _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xfanout46 net48 net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_23_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8732__A2 _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5808_ _1205_ _1197_ _1206_ _0047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6788_ _2096_ _1803_ _2105_ _2106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5546__A2 _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6743__A1 _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8527_ _3051_ _3491_ _3722_ _3498_ _3723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__9048__CLK clknet_leaf_39_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5739_ _1133_ _1151_ _1157_ _0027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8458_ _1645_ _3484_ _3651_ _3461_ _3656_ _3657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__8496__A1 _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7217__C _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7409_ _1586_ _2657_ _2658_ _2659_ _2660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_123_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5849__A3 _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8389_ _1568_ _3588_ _3589_ _3590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_102_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8248__A1 _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8799__A2 _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8420__A1 _2884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6026__A3 _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7223__A2 _2490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8064__B _3294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xwrapped_as2650_62 io_oeb[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_3399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_73 io_oeb[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xwrapped_as2650_84 io_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5785__A2 _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_95 io_oeb[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6734__A1 _2028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7194__I _2464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5707__I _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4611__I _4191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8487__A1 _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7127__C _2398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8487__B2 _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8239__A1 as2650.stack\[7\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6501__A4 _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5442__I _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7462__A2 _4242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7214__A2 _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8411__A1 _2899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5598__B _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7369__I _2561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6273__I _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7760_ _2997_ _2998_ _3003_ _3004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4972_ _0414_ _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6973__A1 _4044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5776__A2 _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6711_ _2029_ _2030_ _2031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7691_ _2891_ _2935_ _2936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8714__A2 _3886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6642_ _4294_ _4301_ _1096_ _1963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_123_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6725__A1 _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5528__A2 _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7922__B1 _3157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8421__C _2687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6573_ _1891_ _1894_ _1895_ _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_34_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8312_ _2403_ _3515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5524_ _0946_ _0960_ _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8243_ net28 _3447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5455_ _0892_ _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__7150__A1 _4049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6876__C _2165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_62_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_62_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_8174_ _3385_ _3398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5386_ _0746_ _0770_ _0824_ _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5700__A2 _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7125_ _2393_ _2396_ _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7056_ _4284_ _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8650__A1 _4195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7453__A2 _4062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8663__I _3835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6007_ _1344_ _1222_ _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4898__S0 _4018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7958_ _2306_ _3178_ _2948_ _3039_ _3195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_43_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6909_ _2207_ _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_126_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7889_ _1797_ _3128_ _3129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8166__B1 _3390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8705__A2 _1859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5519__A2 _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4990__A3 _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8469__A1 _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4742__A3 _4322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7141__A1 _2312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7692__A2 _2931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7995__A3 _3227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5207__A1 _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6093__I _4072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4606__I _4148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5758__A2 _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6955__A1 as2650.r123_2\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_46_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4569__I0 as2650.r123\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9056__D _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5391__B1 _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8748__I _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7652__I _2897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5240_ _0679_ _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4497__A2 _4077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6268__I _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5171_ _0590_ _4378_ _4369_ _0611_ _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_111_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5105__C _4198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5446__A1 _4140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7986__A3 _2393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8930_ _0091_ clknet_leaf_75_wb_clk_i as2650.r123\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput3 io_in[12] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XFILLER_49_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5997__A2 _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8861_ _0022_ clknet_leaf_46_wb_clk_i as2650.stack\[3\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7812_ _3050_ _2987_ _3054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8792_ _0947_ _3940_ _2488_ _2491_ _1288_ _3962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XANTENNA__5749__A2 _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6946__A1 _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7743_ _0723_ _2987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4955_ _0338_ _0341_ _0343_ _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
XANTENNA__8699__A1 _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7674_ as2650.stack\[0\]\[4\] _1193_ _1176_ as2650.stack\[1\]\[4\] _2920_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4886_ _0328_ _0320_ _0325_ _4371_ _0329_ _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6625_ _1891_ _1895_ _1947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_119_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7371__A1 _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6556_ _0837_ _0840_ _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5921__A2 _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5507_ _0944_ _0008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_3_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7123__A1 _4038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6487_ _1809_ _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8226_ _3436_ _3437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6477__A3 _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5438_ _0873_ _0875_ _4291_ _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_133_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8880__CLK clknet_leaf_47_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8157_ _1592_ _3383_ _3384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5082__I _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5369_ _0624_ _0683_ _0686_ _0698_ _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_82_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7108_ _1232_ _0874_ _1235_ _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__6229__A3 _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8623__B2 _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8088_ _1388_ _2494_ _3242_ _3320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_75_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5437__A1 _4163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7039_ _2319_ _2321_ _2322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_142_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4426__I _4006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output15_I net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7362__A1 _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5912__A2 _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7114__A1 _4088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7665__A2 _2285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5676__A1 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6088__I _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7417__A2 _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5428__A1 _4111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8090__A2 _3264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5979__A2 _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_2_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6928__A1 as2650.r123_2\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8252__B _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4740_ _4320_ _4321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4671_ _4226_ _4252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7353__A1 _2439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6410_ _1748_ _1749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__9109__CLK clknet_leaf_9_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7390_ _4364_ _2580_ _2643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6341_ _1648_ _1676_ _1695_ _1697_ _0089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_127_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9060_ _0221_ clknet_leaf_39_wb_clk_i as2650.stack\[6\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6272_ _1638_ _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5667__A1 _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8011_ _2377_ _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5223_ _0562_ _0565_ _0566_ _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__5116__B _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8605__A1 _2862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5154_ as2650.r123\[2\]\[6\] as2650.r123_2\[2\]\[6\] _4013_ _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7408__A2 _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5419__A1 _4302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7959__A3 _3155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5085_ _4002_ _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6092__A1 _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8913_ _0074_ clknet_leaf_9_wb_clk_i as2650.ins_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8844_ _0005_ clknet_leaf_69_wb_clk_i as2650.r123\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6919__A1 _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8775_ _3937_ _3938_ _3946_ _3947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7592__A1 as2650.stack\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5987_ _1373_ _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7726_ _2969_ _2970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4938_ _4324_ _0366_ _0381_ _0002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7344__A1 _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7657_ _2900_ _2865_ _2902_ _2903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__6147__A2 _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4869_ _4178_ _0296_ _0312_ _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6608_ _1928_ _1929_ _1930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7895__A2 _2842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7588_ as2650.stack\[3\]\[3\] _2697_ _1047_ as2650.stack\[2\]\[3\] _2835_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_119_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6539_ _1855_ _1856_ _1861_ _1862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_49_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7647__A2 _2881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8209_ _1684_ _3424_ _3425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8072__A2 _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8056__C _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6083__A1 _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5830__A1 _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_102_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6371__I _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6138__A2 _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7886__A2 _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5897__A1 _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7416__B _2665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7099__B1 _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8247__B _2330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8063__A2 _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6074__A1 _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5821__A1 _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5910_ _1190_ _1301_ _1303_ _0052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6890_ as2650.r123_2\[1\]\[2\] _2193_ _2195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5841_ _1232_ _1235_ _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7574__A1 _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8560_ _3579_ _3752_ _3754_ _3463_ _3517_ _3755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__5585__B1 _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5772_ _1179_ _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4723_ _4303_ _4304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7511_ _2724_ _1278_ _2760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8491_ _3667_ _3669_ _3687_ _3688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7326__A1 _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7442_ _2691_ _2692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4654_ as2650.r123\[1\]\[1\] as2650.r123\[0\]\[1\] as2650.r123_2\[1\]\[1\] as2650.r123_2\[0\]\[1\]
+ as2650.ins_reg\[0\] _4010_ _4235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__9081__CLK clknet_leaf_24_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7373_ _2273_ _2629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8126__I0 _3355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4585_ _4025_ _4166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6324_ _1683_ _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9112_ _0273_ clknet_leaf_47_wb_clk_i as2650.carry vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8826__A1 _2490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9043_ _0204_ clknet_leaf_29_wb_clk_i as2650.pc\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6255_ _1623_ _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6301__A2 _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5206_ _0636_ _0646_ _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6186_ _1560_ _1562_ _1563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_112_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5137_ as2650.r123\[1\]\[4\] _4304_ _0578_ _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8054__A2 _3286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6065__A1 _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7801__A2 _3041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5068_ _0489_ _0509_ _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_83_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4615__A2 _4195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8827_ _3991_ _3992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6191__I _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4704__I _4284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8758_ _2530_ _3282_ _3930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7709_ _2857_ _2939_ _2946_ _2953_ _2954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__7317__A1 _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8689_ _3852_ _0717_ _3865_ _3866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_139_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5879__A1 _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5535__I _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8817__A1 _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4551__A1 _4131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8293__A2 _2749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6366__I _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8045__A2 _4374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5270__I _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5203__C _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7308__A1 _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5445__I _4109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4542__A1 _4119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8808__A1 _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8941__CLK clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6295__A1 _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6040_ _4031_ _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input6_I io_in[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4845__A2 _4412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6276__I _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6047__A1 _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7991_ _2561_ _4262_ _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7795__A1 _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6942_ _2234_ _2235_ _2237_ _0150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7547__A1 _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6873_ _1642_ _2178_ _2182_ _0136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4524__I _4104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8612_ _2306_ _3785_ _3804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_50_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5824_ _1218_ _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8543_ _3055_ _3681_ _3056_ _3739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5755_ _1118_ _1163_ _1168_ _0032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4706_ as2650.halted _4287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8474_ _1412_ _3572_ _3671_ _2622_ _3672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5686_ as2650.pc\[10\] _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7425_ _1417_ _1229_ _2675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4637_ _4217_ _4218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7356_ _2589_ _1054_ _2590_ _2612_ _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4568_ as2650.r123\[0\]\[0\] as2650.r123_2\[0\]\[0\] _4009_ _4149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6307_ _1590_ _1662_ _1669_ _0083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7287_ _2545_ _2546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8275__A2 _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4499_ _4039_ _4080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9026_ _0187_ clknet_leaf_17_wb_clk_i as2650.cycle\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6238_ _1599_ _1604_ _1607_ as2650.stack\[5\]\[0\] _1608_ _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_58_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6169_ _1545_ _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6038__A1 _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6589__A2 _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7011__S _2294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7538__A1 as2650.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4434__I _4014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5974__B _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4772__A1 _4141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8964__CLK clknet_leaf_76_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7710__B2 as2650.stack\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5324__I0 as2650.r123\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5619__A4 _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4609__I _4154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6029__A1 _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8525__B _3493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7777__A1 as2650.pc\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8244__C _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7529__A1 _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6045__B _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5540_ as2650.stack\[4\]\[10\] _0971_ _0973_ as2650.stack\[5\]\[10\] _0976_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_121_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5471_ as2650.psu\[2\] _0891_ _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5307__A3 _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5175__I _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7701__A1 _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7210_ _2345_ _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4515__A1 _4094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4422_ _4002_ _4003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8190_ _3408_ _3409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7141_ _2312_ _4261_ _2331_ _2412_ _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_119_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7072_ _1428_ _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6023_ _1409_ _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5491__A2 _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7974_ as2650.pc\[13\] _1128_ _3139_ _3155_ _3210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_70_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6440__A1 _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5243__A2 _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6925_ _0945_ _1850_ _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_74_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6856_ _2170_ _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout47 net48 net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_126_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5807_ as2650.stack\[1\]\[11\] _1201_ _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7940__A1 _3143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6787_ _0619_ _2056_ _1832_ _2104_ _2105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__8987__CLK clknet_leaf_46_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8526_ _2470_ _3058_ _3721_ _3722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5738_ as2650.stack\[5\]\[12\] _1153_ _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_136_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8457_ _2791_ _2936_ _3655_ _3656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8496__A2 _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5085__I _4002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5669_ _4289_ _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7408_ _1487_ _1586_ _2659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5849__A4 _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8388_ _1631_ _2548_ _2569_ _3589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_117_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8396__I _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6909__I _2207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8248__A2 _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7339_ _2594_ _2595_ _2596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4429__I _4009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9009_ _0170_ clknet_leaf_81_wb_clk_i as2650.r123\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5969__B _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7759__A1 as2650.stack\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6644__I _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8420__A2 _2890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8064__C _3296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6431__A1 _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_63 io_oeb[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_3389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_36_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_as2650_74 io_oeb[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_85 io_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__6982__A2 _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4993__A1 _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8080__B _3270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4745__A1 _4163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7424__B _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8239__A2 _3436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7998__A1 _4364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7998__B2 _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_75_wb_clk_i_I clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5879__B _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7214__A3 _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8411__A2 _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6422__A1 _1629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4971_ _0337_ _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_79_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6973__A2 _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6710_ _2006_ _2009_ _2030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7690_ _2932_ _2934_ _2935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_60_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6641_ _1851_ _1962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7922__A1 _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7922__B2 _2647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6572_ _0335_ _0842_ _1895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8311_ _1502_ _3509_ _3513_ _2625_ _3514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5523_ _4377_ _0947_ _0889_ _0959_ _0929_ _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_121_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6489__A1 _4082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8242_ _1211_ _3438_ _3446_ _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5454_ _0891_ _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7150__A2 _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5385_ _0750_ _0822_ _0823_ _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_8173_ _1675_ _3386_ _3394_ _3397_ _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_114_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7124_ _1429_ _2394_ _2395_ _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_119_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7989__A1 _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7055_ _2334_ _2336_ _1286_ _1223_ _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_115_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8650__A2 _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6006_ _0785_ _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6661__A1 _1942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_31_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_31_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4693__B _4273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_83_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7957_ _1135_ _3193_ _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6908_ _0945_ _2206_ _2207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_70_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7888_ _1255_ _3127_ _3128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8166__A1 _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8166__B2 as2650.stack\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6839_ _1819_ _2152_ _2154_ _2155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7913__A1 _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4712__I _4292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8509_ _3602_ _3705_ _2459_ _3706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8469__A2 _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7141__A2 _4261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8059__C _3243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8641__A2 _3821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6652__A1 _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6404__A1 _1654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5207__A2 _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6955__A2 _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4966__B2 _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8157__A1 _1592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4569__I1 as2650.r123_2\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5391__B2 _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5143__A1 _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6891__A1 _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5170_ _4380_ _0591_ _0610_ _4199_ _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_96_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8632__A2 _3820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5446__A2 _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput4 io_in[13] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_49_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6284__I _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8860_ _0021_ clknet_leaf_47_wb_clk_i as2650.stack\[3\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7811_ _3050_ _3052_ _3053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8791_ _3935_ _3960_ _3961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7742_ _0604_ _0531_ _2986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8148__A1 _2076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4954_ _0396_ _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7329__B _2586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7673_ _0949_ _2918_ _2919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4885_ _4270_ _0301_ _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6624_ as2650.r0\[3\] _0765_ _1946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7371__A2 _2312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6555_ _0834_ _1876_ _1877_ _1878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5506_ _0932_ _0943_ _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_106_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7123__A2 _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6486_ _4098_ _1805_ _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8225_ _3435_ _3436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5437_ _4163_ _4296_ _0874_ _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_82_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7999__B _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8156_ _1173_ _0920_ _3383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5368_ _0802_ _0806_ _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_82_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7107_ _1284_ _2377_ _2378_ _2356_ _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_59_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8623__A2 _3808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5299_ _0652_ _0675_ _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8087_ _3313_ _0428_ _3317_ _3318_ _3319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_60_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5437__A2 _4296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7038_ _1254_ _2320_ _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8387__A1 _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6127__C _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8989_ _0150_ clknet_leaf_67_wb_clk_i as2650.r123_2\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4948__A1 _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8139__A1 _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6143__B _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7362__A2 _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5373__A1 _4179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5373__B2 _4171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8311__A1 _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7114__A2 _4027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5125__A1 _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5273__I _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6873__A1 _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7417__A3 _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5428__A2 _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8252__C _2883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5448__I _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4670_ _4247_ _4250_ _4251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7353__A2 _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6340_ _1696_ _1680_ _1681_ _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6279__I _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6271_ as2650.pc\[4\] _1638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5116__A1 _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5222_ _0661_ _0662_ _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5667__A2 _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8010_ _3244_ _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6864__A1 _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5153_ _0593_ _4021_ _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5911__I _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6616__A1 _1934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5419__A2 _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6467__I1 _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5084_ _0525_ _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8912_ _0073_ clknet_leaf_9_wb_clk_i as2650.ins_reg\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8369__A1 _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8843_ _0004_ clknet_leaf_1_wb_clk_i as2650.r123\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6919__A2 _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7041__A1 _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8774_ _1279_ _3944_ _3945_ _0957_ _3937_ _3946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5986_ _1372_ _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7592__A2 _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7725_ as2650.pc\[6\] _0723_ _2969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4937_ as2650.r123\[1\]\[2\] _4413_ _0380_ _4316_ _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_75_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5358__I _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7656_ _2901_ _2902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4868_ _4168_ _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8541__A1 _3596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7344__A2 _2596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6607_ _1875_ _1901_ _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7587_ _1630_ _2833_ _2834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_20_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4799_ _4249_ _4379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6538_ _1816_ _1857_ _1841_ _1860_ _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_88_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6469_ _1655_ _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_101_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6855__A1 _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8208_ _3411_ _3424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7522__B _2770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8139_ _1580_ _0721_ _3359_ _3367_ _3368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_88_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7280__A1 _4292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5830__A2 _4128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7032__A1 _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8532__A1 _3725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6138__A3 _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7416__C _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7099__A1 _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6099__I as2650.psu\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7099__B2 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5649__A2 _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_106_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8599__A1 net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8247__C _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6449__I1 _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6074__A2 _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5821__A2 _4295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7023__A1 _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5840_ _1233_ _1234_ _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_62_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8870__CLK clknet_leaf_57_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7574__A2 _2816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8771__A1 _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5771_ _1179_ _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5178__I _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7510_ _2739_ _2757_ _2758_ _2759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4722_ _4285_ _4302_ _4137_ _4303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_124_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8490_ _1372_ _0709_ _3687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7326__A2 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7441_ _1045_ _2691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5337__A1 _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4653_ _4212_ _4233_ _4234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__5906__I _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4810__I _4389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7372_ _2624_ _2615_ _2627_ _2628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4584_ _4163_ _4164_ _4165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8126__I1 _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9111_ _0272_ clknet_leaf_41_wb_clk_i as2650.psl\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6323_ as2650.pc\[3\] _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_116_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6837__A1 _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9042_ _0203_ clknet_leaf_29_wb_clk_i as2650.pc\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6254_ _1622_ _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6737__I _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5205_ _0616_ _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6185_ _1561_ _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5136_ _0462_ _0577_ _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7262__A1 _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6065__A2 _4193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5067_ _0410_ _0493_ _0500_ _0508_ _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_38_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8826_ _2490_ _3989_ _3990_ _3991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8762__A1 _3927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8757_ _4308_ _3928_ _2706_ _2646_ _3929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5576__A1 _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5969_ _1039_ _1346_ _1355_ _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_90_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7708_ _1317_ _2433_ _2952_ _2884_ _2953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_55_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8688_ _1040_ _3840_ _3865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8514__A1 _2732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7317__A2 _2450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5328__A1 _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7639_ _1285_ _2884_ _2885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_138_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5879__A2 _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4551__A2 _4059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8817__A2 _2517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6828__A1 _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8893__CLK clknet_leaf_53_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8083__B _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8753__A1 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8811__B _3978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8505__A1 _3515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7308__A2 _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5319__A1 as2650.r0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4542__A2 _4122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8808__A2 _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6819__A1 _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7492__A1 _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5461__I _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6047__A2 _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7244__A1 _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7990_ _1567_ _2417_ _3224_ _3225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_67_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6941_ as2650.r123_2\[0\]\[3\] _2224_ _2236_ _2210_ _2237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_78_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6872_ _1646_ _2179_ _2180_ as2650.stack\[0\]\[5\] _2174_ _2182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__7547__A2 _2794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8611_ _3595_ _3803_ _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5823_ _0860_ _4295_ _0884_ _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_8542_ _3515_ _3736_ _3737_ _3626_ _3738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5754_ as2650.stack\[6\]\[10\] _1166_ _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_56_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_56_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_72_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4705_ _4014_ _4286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8473_ _3667_ _3669_ _3670_ _3671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5685_ _1099_ _1100_ _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4540__I as2650.cycle\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7424_ _4362_ _2672_ _2673_ _2652_ _2674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_124_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4636_ as2650.ins_reg\[0\] as2650.ins_reg\[1\] _4217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_118_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7355_ _2591_ _2609_ _2610_ _2611_ _2334_ _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4567_ as2650.r0\[0\] _4148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6306_ as2650.stack\[4\]\[0\] _1665_ _1668_ _1661_ _1669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_104_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7286_ _2415_ _2545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4498_ _4072_ _4078_ _4079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9025_ _0186_ clknet_3_3_0_wb_clk_i as2650.halted vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6237_ _1593_ _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6168_ _4073_ _1070_ _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7800__B _2789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5119_ _0560_ _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6099_ as2650.psu\[3\] _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_85_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_26_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_3_3_0_wb_clk_i clknet_0_wb_clk_i clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__7538__A2 _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8809_ _1258_ _1260_ _1263_ _3976_ _3977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_41_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5021__I0 as2650.r123\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5721__A1 _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5324__I1 as2650.r123_2\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_65_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6029__A2 _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5237__B1 _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7777__A2 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9071__CLK clknet_leaf_42_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4625__I as2650.psl\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7529__A2 _2776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6045__C _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7157__B _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5960__A1 _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4763__A2 _4298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5470_ _0907_ _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_117_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7701__A2 _2868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5307__A4 _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4421_ _4001_ _4002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4515__A2 _4095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5712__A1 _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5712__B2 as2650.r123_2\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7140_ _2407_ _2411_ _2412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7465__A1 _1597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7071_ _1252_ _1544_ _2352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_59_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6022_ _0540_ _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_95_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5779__A1 _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7973_ _2462_ _3208_ _3209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6924_ _0959_ _2213_ _2221_ _2222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6440__A2 _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6855_ _1713_ _0977_ _1750_ _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8451__B _3649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout48 net49 net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_11_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5806_ _1125_ _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6786_ _1808_ _2102_ _2103_ _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7940__A2 _3145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8525_ _3326_ _3719_ _3493_ _3720_ _3721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5737_ _1126_ _1150_ _1156_ _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8456_ _1644_ _3480_ _3653_ _3654_ _3655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5668_ _1097_ _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_129_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7407_ _1500_ _2354_ _1370_ _2658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_136_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4619_ _4199_ _4200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8387_ _1256_ _2701_ _3587_ _3588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5599_ as2650.stack\[0\]\[14\] _0953_ _0907_ as2650.stack\[1\]\[14\] _1031_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_117_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7338_ _4121_ _4103_ _2595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7514__C _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7456__A1 _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7269_ _0799_ _2503_ _2529_ _0185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9008_ _0169_ clknet_leaf_76_wb_clk_i as2650.r123\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9094__CLK clknet_leaf_51_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8405__B1 _3540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4690__A1 _4265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7759__A2 _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output38_I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5234__A3 _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6431__A2 _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_64 io_oeb[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4442__A1 _4017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_75 io_oeb[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8708__A1 _3880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_as2650_86 io_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_109_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8931__CLK clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8184__A2 _3390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6195__A1 _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7931__A2 _3147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5276__I _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5942__A1 _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4745__A2 _4145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7695__A1 _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_1_wb_clk_i clknet_3_0_0_wb_clk_i clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_108_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7424__C _2652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5170__A2 _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7998__A2 _4060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5879__C _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4681__A1 _4093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4970_ _0412_ _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_63_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6973__A3 _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5895__B _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8175__A2 _3393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6640_ _1852_ _1923_ _1924_ _1961_ _0124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6186__A1 _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7922__A2 _3150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6571_ _0416_ _0560_ _1894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5933__A1 _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8310_ _3468_ _3512_ _3513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5522_ _0951_ _0955_ _0956_ _0958_ _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_121_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8241_ as2650.stack\[7\]\[14\] _3436_ _3446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6489__A2 _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5453_ _0890_ as2650.psu\[1\] _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7150__A3 _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8172_ _1679_ _3395_ _3396_ _3397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5384_ _0755_ _0821_ _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_114_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7123_ _4038_ _1543_ _2289_ _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_119_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7989__A2 _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7054_ _2335_ _2336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7350__B _2595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6005_ _1363_ _1384_ _1391_ _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_86_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4672__A1 _4243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8954__CLK clknet_leaf_47_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_71_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_71_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_7956_ _1128_ _3139_ _3141_ _3193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6907_ _4086_ _1806_ _2205_ _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7887_ _0349_ _2260_ _3126_ _3127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7576__I _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6480__I _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6177__A1 _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6838_ _0787_ _1855_ _2153_ _1821_ _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7913__A2 _2593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5924__A1 _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5096__I net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6769_ _1937_ _2087_ _2088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8508_ _3020_ _3704_ _3705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7677__A1 _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8439_ _1282_ _3565_ _2287_ _3637_ _3638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__5824__I _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7429__A1 _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8356__B _2485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6652__A2 _4116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6404__A2 _1712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7486__I _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8157__A2 _3383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4903__I net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6168__A1 _4073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7668__A1 _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8110__I _2626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6340__A1 _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5143__A2 _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6891__A2 _2071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8977__CLK clknet_leaf_58_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7840__A1 _3051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xinput5 io_in[5] net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7810_ _1793_ _3010_ _3052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_64_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8790_ _1559_ _3920_ _3960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_92_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7741_ _1650_ _2984_ _2985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4953_ _4115_ _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8148__A2 _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4813__I _4392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7672_ as2650.stack\[3\]\[4\] _1663_ _2918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4884_ as2650.addr_buff\[6\] _4266_ _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6623_ _1941_ _1944_ _1945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7371__A3 _4074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6554_ _0836_ _0852_ _1877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_118_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5382__A2 _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7659__A1 _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5505_ _0933_ _0942_ _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5644__I _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6485_ _1807_ _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7123__A3 _2289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8224_ _1145_ _3383_ _3435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5436_ _4067_ _4144_ _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5134__A2 _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6331__A1 _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_3_1_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8155_ _1653_ _3245_ _3382_ _2730_ _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5367_ _0682_ _0684_ _0805_ _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7106_ _4307_ _1436_ _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8086_ _3303_ _2014_ _1385_ _3318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_99_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5298_ _0702_ _0737_ _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7037_ _1845_ _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7831__A1 _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5437__A3 _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4645__A1 _4225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8387__A2 _2701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6398__A1 _1738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_8988_ _0149_ clknet_leaf_69_wb_clk_i as2650.r123_2\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7939_ _2882_ _3176_ _2894_ _3177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5819__I _4307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8139__A2 _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6143__C _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7898__A1 _2831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7362__A3 _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6570__A1 _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4879__B _4153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7255__B _2518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7114__A3 _4400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5125__A2 _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6322__A1 _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8075__A1 _3297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8086__B _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7822__A1 _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5503__B _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5428__A3 _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6385__I _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4636__A1 as2650.ins_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8814__B _3974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6389__A1 _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7050__A2 _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4939__A2 _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5061__A1 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4633__I _4213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7889__A1 _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7353__A3 _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5116__A2 _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6270_ _1594_ _1637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6313__A1 _1611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5221_ _0533_ _4318_ _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__9005__CLK clknet_leaf_76_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8066__A1 _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5152_ _0592_ _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6616__A2 _1937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5083_ _0524_ _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8911_ _0072_ clknet_leaf_10_wb_clk_i as2650.ins_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8842_ _0003_ clknet_leaf_1_wb_clk_i as2650.r123\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7041__A2 _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8773_ _0965_ _1279_ _3945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5985_ _1371_ _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5639__I _4080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5052__A1 as2650.holding_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7724_ _1738_ _2967_ _2968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4936_ _0378_ _0379_ _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_40_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7655_ net9 _0420_ _2901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_21_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4867_ _4171_ _0303_ _0310_ _4348_ _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_123_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6606_ _1878_ _1900_ _1928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7586_ as2650.pc\[2\] as2650.pc\[1\] as2650.pc\[0\] _2833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_4798_ _4198_ _4378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6537_ _1859_ _1813_ _1860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6468_ _1792_ _0121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8207_ _1675_ _3410_ _3422_ _3423_ _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_133_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5419_ _4302_ _0857_ _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6855__A2 _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6399_ as2650.stack\[3\]\[6\] _1731_ _1739_ _1710_ _1740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_121_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4866__A1 _4335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8057__A1 _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4866__B2 _4343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8138_ _1386_ _3263_ _3259_ _3366_ _3264_ _0726_ _3367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_134_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7804__A1 _2438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4718__I _4298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8069_ _0370_ _3246_ _3301_ _1527_ _3302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_82_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7280__A2 _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5291__A1 _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8126__S _3244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5830__A3 _4145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7032__A2 _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5043__A1 _4324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4453__I _4033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5594__A2 _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5993__B _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9028__CLK clknet_leaf_17_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8296__A1 _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7099__A2 _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8809__B _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4628__I _4208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6074__A3 _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5821__A3 _4312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7023__A2 _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8220__A1 _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_opt_1_0_wb_clk_i_I clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5034__A1 _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8771__A2 _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_50_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5770_ _1178_ _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5585__A2 _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6782__A1 _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4721_ _4290_ _4294_ _4301_ _4302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_72_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7440_ _2316_ _2690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4652_ as2650.r123\[2\]\[1\] as2650.r123_2\[2\]\[1\] _4010_ _4233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6534__A1 _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7371_ _1231_ _2312_ _4074_ _2626_ _2627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_50_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4583_ _4071_ _4164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_9110_ _0271_ clknet_leaf_9_wb_clk_i as2650.ins_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6322_ _1675_ _1676_ _1678_ _1682_ _0085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_115_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7623__B _2869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9041_ _0202_ clknet_leaf_31_wb_clk_i as2650.pc\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6253_ _1621_ _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4848__A1 _4289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8039__A1 _3271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5204_ _0632_ _0635_ _0644_ _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_69_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6184_ _4032_ _1427_ _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4538__I as2650.cycle\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5135_ _0479_ _0575_ _0576_ _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7798__B1 _3037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7262__A2 _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6065__A3 _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5066_ _4179_ _0503_ _0507_ _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8211__A1 _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8825_ _1542_ _4311_ _3975_ _3990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__5025__A1 _4375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6773__A1 _2028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8756_ _4314_ _3251_ _3928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5968_ _1354_ _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7707_ _2446_ _2931_ _2951_ _2952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4919_ _4258_ _0331_ _0362_ _4367_ _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_8687_ _3851_ _3863_ _3864_ _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7584__I _2438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6702__B _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5899_ _1293_ _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7638_ _2883_ _2884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6525__A1 _1847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7517__C _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7569_ as2650.stack\[3\]\[2\] _1297_ _1176_ as2650.stack\[1\]\[2\] _2817_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_140_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8278__B2 _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_55_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5264__A1 _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5016__A1 _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8753__A2 _2676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5567__A2 _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6764__A1 _4209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7708__B _2884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8505__A2 _3698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7713__B1 _2956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8269__A1 _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7492__A2 _4233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7244__A2 _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5255__A1 _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6940_ _2023_ _2024_ _2208_ _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_81_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6871_ _2177_ _2178_ _2181_ _0135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5007__A1 _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8744__A2 _3914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8610_ net39 _3523_ _3802_ _3803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_90_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5822_ _1216_ _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6755__A1 _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5558__A2 _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8541_ _3596_ _3719_ _3737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7618__B _2864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5753_ _1110_ _1163_ _1167_ _0031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4704_ _4284_ _4285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8472_ _3667_ _3669_ _3468_ _3670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6507__A1 _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5684_ _1087_ _1110_ _1112_ _0017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_136_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7423_ _1342_ _1063_ _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_135_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4635_ _4214_ _4215_ _4216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7180__A1 _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7354_ _2410_ _2611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_25_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_25_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_85_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4566_ _4146_ _4147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5730__A2 _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7353__B _2596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6305_ _1667_ _1665_ _1668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7285_ _2434_ _2539_ _2540_ _2541_ _2543_ _2544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_103_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4497_ _4073_ _4077_ _4078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_9024_ _0185_ clknet_leaf_7_wb_clk_i as2650.holding_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6236_ _1606_ _1607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5494__A1 _4283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6167_ _1543_ _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_112_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8432__A1 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5118_ as2650.r123\[0\]\[4\] as2650.r123_2\[0\]\[4\] as2650.psl\[4\] _0560_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_3506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6098_ _0430_ _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_3517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5246__A1 _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6483__I _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5049_ _0419_ _0421_ _0423_ _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_72_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6994__A1 _4105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5797__A2 _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8735__A2 _3906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8808_ _1560_ _1500_ _3976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6746__A1 _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8739_ _3911_ _2488_ _3303_ _3912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_41_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8499__A1 _3603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7171__A1 _2436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5021__I1 as2650.r123_2\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8860__CLK clknet_leaf_47_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8423__A1 _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8094__B _3324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5237__A1 as2650.r123\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5237__B2 _4316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6985__A1 _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6326__C _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8822__B as2650.psl\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8187__B1 _3390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8726__A2 _3893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4641__I _4221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5960__A2 _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4420_ as2650.ins_reg\[0\] _4001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7465__A2 _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7070_ _2344_ _2348_ _2350_ _2351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8662__A1 _3838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6021_ _1399_ _1401_ _1405_ _1407_ _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA_clkbuf_3_6_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7217__A2 _2484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5228__A1 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7399__I _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5779__A2 _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7972_ as2650.pc\[14\] _3207_ _3208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_54_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6923_ _2214_ _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8717__A2 _2096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6728__A1 _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6854_ _2168_ _2169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7925__B1 _3157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8451__C _2580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout49 net50 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5805_ _1203_ _1197_ _1204_ _0046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_56_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6785_ _0587_ _1966_ _2103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8023__I _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8524_ _2252_ _3326_ _3720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5736_ as2650.stack\[5\]\[11\] _1153_ _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5951__A2 _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7153__A1 _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8455_ _2668_ _3654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5667_ _1094_ _1096_ _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4618_ _4198_ _4199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7406_ _2656_ _1370_ _2657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8386_ _2852_ _3586_ _3587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8883__CLK clknet_leaf_51_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6900__A1 _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5598_ as2650.stack\[7\]\[14\] _0977_ _0957_ _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7337_ _2593_ _2594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6478__I _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4549_ _4128_ _4129_ _4130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7456__A2 _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7268_ _2503_ _2528_ _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9007_ _0168_ clknet_leaf_76_wb_clk_i as2650.r123\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6219_ _1589_ _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7199_ _2469_ _2470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_63_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8405__A1 _2899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5219__A1 _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4690__A2 _4270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4726__I _4291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6967__A1 _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_65 io_oeb[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_76 io_oeb[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_87 io_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6195__A2 _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7695__A2 _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8817__B _3978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7721__B _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7998__A3 _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4681__A2 _4096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6958__A1 as2650.r123_2\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6851__I _2165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7383__A1 _2613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6186__A2 _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6570_ _0762_ _1891_ _1892_ _0848_ _1893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_32_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5933__A2 _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5521_ as2650.stack\[7\]\[9\] _0893_ _0952_ as2650.stack\[6\]\[9\] _0957_ _0958_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7135__A1 _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8240_ _1209_ _3438_ _3445_ _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5452_ as2650.psu\[0\] _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6298__I _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8171_ _3384_ _3396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5383_ _0755_ _0821_ _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7122_ _1342_ _2277_ _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7053_ _1272_ _2335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7989__A3 _2656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5930__I _4293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6004_ _1385_ _0782_ _1390_ _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_101_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6949__A1 _2106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7955_ _2830_ _3190_ _3192_ _0208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_70_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5621__A1 _4288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6906_ _1842_ _1911_ _1829_ _1802_ _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_7886_ as2650.addr_buff\[2\] _0290_ _3126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6837_ _1519_ _1854_ _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6177__A2 _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7374__A1 _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6768_ _2081_ _2086_ _2087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5924__A2 _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_40_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_40_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_104_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8507_ _3021_ _3703_ _3704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5719_ _1142_ _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7126__A1 _4108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6699_ _0414_ _1973_ _2019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8438_ _3634_ _3635_ _3636_ _3637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9061__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8369_ _1406_ _3565_ _3464_ _3569_ _3570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_123_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6001__I _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7429__A2 _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6652__A3 _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4663__A2 _4106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7601__A2 _2786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5073__C1 _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8091__C _2639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7365__A1 _2439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6168__A2 _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5915__A2 _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7117__A1 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5679__A1 _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7840__A2 _2686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5851__A1 _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput6 io_in[6] net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5603__A1 _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5603__B2 _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7740_ _1643_ _1638_ _2907_ _2984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4952_ as2650.holding_reg\[3\] _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_45_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4883_ _0321_ _0326_ _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7671_ as2650.stack\[6\]\[4\] _2692_ _2695_ as2650.stack\[5\]\[4\] _2917_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_6622_ _1942_ _1943_ _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_14_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9084__CLK clknet_leaf_25_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6553_ _0836_ _0852_ _1876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7108__A1 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5504_ _0941_ _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7659__A2 _2593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6484_ _4366_ _1806_ _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5435_ _0504_ _4299_ _4300_ _0872_ _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_8223_ _1698_ _3419_ _3434_ _0234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_127_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8608__A1 _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5366_ _0698_ _0691_ _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8154_ _3372_ _3381_ _3276_ _3382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7105_ _0934_ _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8085_ _0470_ _3246_ _3316_ _1528_ _3317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__8084__A2 _2841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5297_ _0293_ _0732_ _0736_ _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_82_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8921__CLK clknet_leaf_33_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7036_ _2318_ _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7831__A2 _3053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5842__A1 _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8987_ _0148_ clknet_leaf_46_wb_clk_i as2650.r123_2\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8792__B1 _2491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7938_ _2885_ _3168_ _3175_ _2758_ _3176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_43_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7347__A1 _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7869_ _3083_ _2686_ _3109_ _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_109_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5835__I _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4581__A1 as2650.holding_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_2_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6086__A1 _1470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5503__C _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7822__A2 _4215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5833__A1 _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4636__A2 as2650.ins_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8814__C _3981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7586__A1 as2650.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5597__B1 _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5597__C2 _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5061__A2 _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7338__A1 _4121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6010__A1 _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6561__A2 _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8302__A3 _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6849__B1 _2163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8944__CLK clknet_leaf_56_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6313__A2 _1662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5220_ _0565_ _0660_ _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_124_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5521__B1 _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4875__A2 _4232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5151_ as2650.r0\[6\] _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5480__I _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5082_ _0523_ _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8910_ _0071_ clknet_leaf_9_wb_clk_i as2650.ins_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8841_ _0002_ clknet_leaf_2_wb_clk_i as2650.r123\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_112_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8772_ _3942_ _3943_ _3944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5984_ _0723_ _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5052__A2 _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7723_ _1644_ _2930_ _2967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4935_ _0376_ _0377_ _0284_ _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_36_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7654_ _2899_ _0340_ _2900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4866_ _4335_ _0307_ _0309_ _4343_ _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7356__B _2590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6605_ _1869_ _1925_ _1926_ _1927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7585_ _2824_ _2832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4797_ _4376_ _4377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4563__A1 _4026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6536_ _1858_ _1859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7501__A1 _4393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6467_ _1791_ _1028_ _1778_ _1792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_133_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8206_ _1624_ _3416_ _3417_ _3423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5418_ _0820_ _0856_ _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA_clkbuf_leaf_45_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6855__A3 _1750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6398_ _1738_ _1714_ _1739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_47_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8137_ _1381_ _0646_ _3364_ _1422_ _3365_ _3366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5349_ _4246_ _0787_ _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8057__A2 _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8068_ _3298_ _3299_ _0935_ _3300_ _3301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_102_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7019_ as2650.addr_buff\[4\] _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_56_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7568__A1 as2650.stack\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5043__A2 _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8650__B _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5993__C _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8097__B _3270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6396__I as2650.pc\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5514__B _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6059__A1 _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5282__A2 _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8220__A2 _3419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7020__I _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4720_ _4296_ _4299_ _4300_ _4301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4651_ _4230_ _4231_ _4232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__6534__A2 _1843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4545__A1 _4064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7370_ _2625_ _2626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4582_ _4140_ _4163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_116_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6321_ _1679_ _1680_ _1681_ _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6252_ as2650.pc\[2\] _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9040_ _0201_ clknet_leaf_31_wb_clk_i as2650.pc\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4848__A2 _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5203_ _0312_ _0639_ _0643_ _0403_ _0299_ _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_115_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6183_ _1057_ _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_131_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8039__A2 _4279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5134_ _0479_ _0574_ _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7798__A1 _3029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7798__B2 _3039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5065_ _4168_ _0488_ _0506_ _4299_ _4165_ _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_38_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8824_ _1261_ _1221_ _3249_ _3989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8211__A2 _3419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6222__A1 _1592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8755_ _2257_ _3926_ _3927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5967_ _1353_ _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7706_ _2947_ _2935_ _2950_ _2951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4918_ _0334_ _4199_ _4257_ _0361_ _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_8686_ net20 _3839_ _3864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5898_ _0940_ _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7637_ _2417_ _2883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4849_ _0292_ _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6525__A2 _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4536__A1 _4109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7568_ as2650.stack\[2\]\[2\] _2691_ _1193_ as2650.stack\[0\]\[2\] _2816_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_105_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_1_wb_clk_i_I clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6519_ _1814_ _1842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7499_ as2650.pc\[1\] net6 _2748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_106_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9169_ net47 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7105__I _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7789__A1 _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8450__A2 _3648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8202__A2 _3412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5016__A2 _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8380__B _3580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7961__A1 _4095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6764__A2 _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5295__I _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7713__B2 as2650.stack\[5\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8269__A2 _2489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7015__I _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6854__I _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8441__A2 _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6452__A1 as2650.stack\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6870_ _1639_ _2179_ _2180_ as2650.stack\[0\]\[4\] _2174_ _2181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__6204__A1 _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5821_ _0860_ _4295_ _4312_ _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7952__A1 _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7952__B2 _2688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8540_ _3340_ _3729_ _3735_ _3507_ _3736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4766__A1 _4344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5752_ as2650.stack\[6\]\[9\] _1166_ _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7004__I0 _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4703_ net10 _4284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_8471_ _3640_ _3644_ _3668_ _3669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_30_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7704__A1 _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5683_ as2650.stack\[3\]\[9\] _1111_ _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_72_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7422_ _1065_ _2325_ _1071_ _2672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4634_ as2650.r123\[2\]\[7\] as2650.r123_2\[2\]\[7\] _4013_ _4215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7180__A2 _4089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7353_ _2439_ _1346_ _1452_ _2596_ _2610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__5191__A1 _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4565_ _4142_ _4145_ _4146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8449__C _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6304_ _1666_ _1667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7284_ _2434_ _2542_ _2543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4496_ _4076_ _4077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9023_ _0184_ clknet_3_2_0_wb_clk_i as2650.holding_reg\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6235_ _1044_ _0971_ _1605_ _1606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
Xclkbuf_leaf_65_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_65_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6691__A1 _1962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6166_ _1427_ _4054_ _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_98_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5117_ _0463_ _0478_ _0480_ _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6097_ _4006_ _1482_ _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5246__A2 _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5048_ as2650.holding_reg\[4\] _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9018__CLK clknet_leaf_7_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6994__A2 _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8196__A1 _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8807_ _1553_ _1370_ _2530_ _2548_ _3975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_80_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7595__I _2690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6999_ _2285_ _2287_ _2289_ _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8738_ _1266_ _3911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_41_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6432__C _1744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8669_ _3836_ _3849_ _3850_ _0264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7171__A2 _2442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7544__B _2791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5182__A1 as2650.holding_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7459__B1 _2285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8120__A1 _3344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4459__I _4039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5237__A2 _4413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6985__A2 _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8187__A1 _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7234__I0 as2650.holding_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7719__B _2791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5960__A3 _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4920__A1 _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8111__A1 _3340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6122__B1 _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8662__A2 _3258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6673__A1 _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6020_ _1406_ _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_136_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input4_I io_in[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8414__A2 _3613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5228__A2 _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7971_ as2650.pc\[13\] as2650.pc\[12\] _1120_ _3140_ _3207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6922_ _1777_ _2219_ _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_130_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6853_ _1747_ _1298_ _1601_ _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__7925__A1 _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7925__B2 _2689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5804_ as2650.stack\[1\]\[10\] _1201_ _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6784_ _1022_ _1908_ _1829_ _2101_ _2102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_8523_ _3716_ _3718_ _3719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_50_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5735_ _1118_ _1150_ _1155_ _0025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8454_ _2949_ _3652_ _3653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5666_ _1095_ _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8350__A1 _3549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7405_ _4131_ _2656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_129_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4617_ _4196_ _4197_ _4198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8385_ _2897_ _3564_ _3586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6900__A2 _2192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5597_ as2650.stack\[6\]\[14\] _0952_ _0988_ as2650.stack\[4\]\[14\] as2650.stack\[5\]\[14\]
+ _0908_ _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_89_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7336_ _2320_ _2593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4548_ _4115_ _4129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8102__A1 _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7267_ _1523_ _2517_ _1526_ _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4479_ _4059_ _4060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_9006_ _0167_ clknet_leaf_77_wb_clk_i as2650.r123\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6218_ _1588_ _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7198_ _2417_ _2469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8405__A2 _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6149_ as2650.r123_2\[3\]\[0\] _1534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5219__A2 _4414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6416__A1 _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6416__B2 as2650.stack\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6967__A2 _2257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4978__A1 _4213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_55 io_oeb[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_66 io_oeb[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_77 io_oeb[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_54_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_88 io_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7274__B _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5155__A1 _4214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8644__A2 _3819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6655__A1 _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6958__A2 _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4969__A1 _4147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7907__A1 _3143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5748__I _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5520_ _0923_ _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_125_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7135__A2 _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5451_ _4290_ _0888_ _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8170_ _3387_ _3395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5382_ _0747_ _0761_ _0768_ _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_7121_ _4364_ _2290_ _2393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8635__A2 _3820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6646__A1 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7052_ _1251_ _2334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6003_ _0428_ _0714_ _1386_ _1389_ _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_45_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7071__A1 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7954_ _1130_ _2829_ _3191_ _3192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5621__A2 _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6905_ _2163_ _2186_ _2204_ _0146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7885_ _3120_ _3124_ _3125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_51_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8034__I _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7078__C _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6836_ _4225_ _0782_ _1813_ _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8571__A1 _3725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7374__A2 _2629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8850__CLK clknet_leaf_67_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6767_ _2084_ _2085_ _2086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7873__I _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8506_ _2970_ _3681_ _3703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5718_ as2650.r123\[0\]\[6\] _1113_ _1141_ _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6698_ _2014_ _1839_ _2017_ _1816_ _2018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7126__A2 _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5137__A1 as2650.r123\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8437_ _3634_ _3635_ _4060_ _3636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5649_ _1074_ _1078_ _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_108_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_80_wb_clk_i clknet_3_0_0_wb_clk_i clknet_leaf_80_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_139_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8368_ _3565_ _3568_ _3569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_123_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7319_ _1257_ _2576_ _2440_ _2574_ _2577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_105_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8087__B1 _3317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8299_ _1496_ _4278_ _3502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_2_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4737__I _4149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5073__C2 _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4472__I as2650.cycle\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8562__A1 _2862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7365__A2 _2620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5376__A1 _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7117__A2 _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6876__A1 _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput7 io_in[7] net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8282__C _3485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8873__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5603__A2 _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4951_ _0384_ _0393_ _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5478__I _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7670_ as2650.stack\[7\]\[4\] _2697_ _2836_ as2650.stack\[4\]\[4\] _2916_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4882_ _0322_ _4389_ _0325_ _4356_ _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_4
XFILLER_71_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7356__A2 _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8553__A1 _3062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6621_ _4382_ _1935_ _0467_ _0592_ _1943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5367__A1 _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6552_ _0758_ _0837_ _0831_ _1874_ _1875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__8305__A1 _3465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7108__A2 _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5503_ _4290_ _0939_ _0869_ _0940_ _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_119_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6483_ _1805_ _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6102__I _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8222_ as2650.stack\[7\]\[7\] _3424_ _3433_ _3408_ _3434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5434_ _4004_ _0521_ _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_105_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_35_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8153_ _1569_ _0787_ _1397_ _3380_ _2651_ _1340_ _3381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__8608__A2 _3483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5365_ _0622_ _0803_ _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6619__A1 _4208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7104_ _4049_ _1561_ _2376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_141_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8084_ _3253_ _2841_ _3314_ _3315_ _0935_ _3316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_5296_ _4280_ _0735_ _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4557__I _4137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7292__A1 _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7035_ _1344_ _1460_ _2318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8029__I _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8986_ _0147_ clknet_leaf_69_wb_clk_i as2650.r123_2\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8792__A1 _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8792__B2 _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7937_ _2788_ _3174_ _3175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7868_ _2685_ _3108_ _2927_ _3109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7347__A2 _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6819_ _0680_ _0720_ _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7799_ _2892_ _3024_ _3042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_clkbuf_leaf_74_wb_clk_i_I clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6858__A1 _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6012__I _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5530__A1 _4017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5833__A2 _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8896__CLK clknet_leaf_51_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7035__A1 _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7586__A2 as2650.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8783__A1 _1610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7338__A2 _4103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6010__A2 _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8402__I _2559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7446__C _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6849__A1 _2013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6849__B2 _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5521__B2 as2650.stack\[6\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5150_ _0492_ _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7274__A1 _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5081_ as2650.r123\[0\]\[5\] as2650.r123_2\[0\]\[5\] as2650.psl\[4\] _0523_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_57_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8840_ _0001_ clknet_leaf_70_wb_clk_i as2650.r123\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7577__A2 _2777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8774__A1 _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8774__B2 _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8771_ _1575_ _1288_ _1336_ _3943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__9051__CLK clknet_leaf_66_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5983_ _1369_ _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7722_ _2929_ _2966_ _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4934_ _0284_ _0376_ _0377_ _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_52_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8526__A1 _2470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8740__C _3313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7653_ _0429_ _2899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_4865_ _0298_ _0308_ _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_123_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6604_ _1873_ _1902_ _1926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7356__C _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7584_ _2438_ _2831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4796_ _4375_ _4376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6535_ _1069_ _1269_ _1858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4563__A2 _4143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6466_ _1738_ _1782_ _1790_ _1791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7501__A2 _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7372__B _2627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8205_ as2650.stack\[7\]\[2\] _3413_ _3422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5417_ _0825_ _0855_ _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6397_ _1737_ _1738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8136_ _1479_ _4223_ _3365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5348_ _4221_ _0786_ _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_88_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8067_ _0879_ _2822_ _3300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5279_ _4394_ _0615_ _0580_ _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_130_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7018_ _2301_ _2302_ _2305_ _0158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7017__A1 _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5028__B1 _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7568__A2 _2691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8969_ _0130_ clknet_leaf_4_wb_clk_i as2650.r123_2\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5503__A1 _4290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6059__A2 _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9074__CLK clknet_leaf_51_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4490__A1 _4026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8756__A1 _4314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5990__A1 _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4793__A2 _4332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4660__I net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4650_ _4001_ as2650.ins_reg\[1\] _4231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6534__A3 _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput10 wb_rst_i net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyd_1
XANTENNA__4545__A2 _4026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4581_ as2650.holding_reg\[0\] _4161_ _4162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6320_ _1660_ _1681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_122_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7495__A1 _2594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7192__B _2456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6251_ _1619_ _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5202_ _0640_ _0537_ _0642_ _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6182_ _1399_ _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5133_ _0559_ _0574_ _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_69_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7798__A2 _3031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5064_ _4193_ _0427_ _0505_ _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_42_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4835__I _4414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7211__I _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8747__A1 _3910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8823_ _3978_ _3987_ _3988_ _3659_ _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_92_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5025__A3 _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6222__A2 _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8754_ _2542_ _2325_ _2598_ _3926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_53_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5966_ _1352_ _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7705_ _1440_ _2948_ _2949_ _2950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4917_ _4240_ _4239_ _0360_ _4198_ _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5981__A1 _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8685_ _3852_ _0681_ _3862_ _3863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5666__I _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5897_ _1279_ _1291_ _1277_ _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8042__I _3243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7636_ _2707_ _2882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7183__B1 _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4848_ _4289_ _0291_ _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7722__A2 _2966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7567_ _2592_ _2814_ _2815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5733__A1 _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4536__A2 _4112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4779_ _4358_ _4359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6518_ _1840_ _1806_ _1841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7498_ _1335_ _2737_ _2734_ _2747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_49_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6449_ _1776_ _1777_ _1778_ _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9168_ net47 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9097__CLK clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7238__A1 _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8119_ _0526_ _2377_ _3348_ _1527_ _3349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_103_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9099_ _0260_ clknet_leaf_50_wb_clk_i as2650.stack\[4\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7789__A2 _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8934__CLK clknet_opt_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7410__A1 _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8380__C _2629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7961__A2 _2861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7713__A2 _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5724__A1 _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6200__I _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8836__B as2650.psu\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7229__A1 _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6452__A2 _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8729__A1 _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8729__B2 _2096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8571__B _4092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7401__A1 _4261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6204__A2 _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5820_ _4314_ _0926_ _0885_ _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_23_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5751_ _1161_ _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5963__A1 _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6091__B _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7004__I1 _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4702_ _4139_ _4186_ _4282_ _4283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_72_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8470_ _3641_ _3668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_124_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5682_ _1085_ _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7704__A2 _2860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7421_ _2396_ _2454_ _2667_ _2670_ _2671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_72_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4633_ _4213_ _4214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5715__A1 _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7180__A3 _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7352_ _2336_ _2602_ _2604_ _2608_ _2609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_102_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4564_ _4144_ _4145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7468__A1 _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6303_ _1596_ _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7283_ _1065_ _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4495_ _4041_ _4075_ _4076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5479__B1 _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6110__I net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9022_ _0183_ clknet_leaf_7_wb_clk_i as2650.holding_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6234_ _1082_ _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6140__A1 _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8746__B _2534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8417__B1 _3601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6691__A2 _1979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6165_ _4006_ _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5116_ _0293_ _0511_ _0557_ _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_69_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6096_ _1224_ _1417_ _4128_ _4335_ _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_131_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8957__CLK clknet_leaf_56_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5047_ _0486_ _0488_ _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_34_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_34_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_38_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8196__A2 _3383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8806_ _1258_ _1416_ _3974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6998_ _2288_ _2272_ _2289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7943__A2 _3180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8737_ _3904_ _3908_ _3909_ _3869_ _3910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_94_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5949_ _1335_ _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8668_ net43 _3846_ _3850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_16_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7619_ _2863_ _2810_ _2864_ _2866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__5706__A1 _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8599_ net39 _3791_ _3792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5706__B2 as2650.r123_2\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5182__A2 _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7459__A1 _4243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7459__B2 as2650.addr_buff\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6020__I _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6131__A1 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6131__B2 _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4693__A1 _4264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5080__B _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4475__I _4055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8391__B _3591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7786__I _2704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4996__A2 _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7234__I1 _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6198__A1 _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9112__CLK clknet_leaf_47_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4748__A2 _4238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_73_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7698__A1 _2940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4920__A2 _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8111__A2 _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6122__A1 _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7870__A1 _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6673__A2 _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7970_ _3205_ _3206_ _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4436__A1 _4015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6921_ _2218_ _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8178__A2 _3393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6852_ _2166_ _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6189__A1 _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7925__A2 _2690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5803_ _1117_ _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6783_ _1971_ _2100_ _2101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8522_ _3717_ _3699_ _3718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5734_ as2650.stack\[5\]\[10\] _1153_ _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_17_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8453_ _2868_ _3631_ _3652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5665_ _4015_ _4288_ _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8320__I _3459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7404_ _2589_ _4048_ _2590_ _2655_ _0194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_50_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4616_ _4082_ _4112_ _4197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8384_ _2788_ _2849_ _3585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5596_ _0711_ _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7335_ _2464_ _2592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4547_ _4087_ _4128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8102__A2 _3331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7266_ _2527_ _0184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4478_ _4057_ _4058_ _4059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7380__B _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9005_ _0166_ clknet_leaf_76_wb_clk_i as2650.r123\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7861__A1 _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6217_ _4188_ _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_132_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7197_ _1066_ _2465_ _2456_ _2467_ _2468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_48_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6148_ _1468_ _1532_ _1533_ _1295_ _0060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_46_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6079_ _0640_ _1462_ _1464_ _1254_ _1465_ _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XTAP_3327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4978__A2 _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_as2650_56 io_oeb[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8169__A2 _3393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_67 io_oeb[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_78 io_oeb[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_89 io_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5927__A1 _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6015__I net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5854__I _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8230__I _3435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5155__A2 _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7852__A1 _2788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7449__C _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7907__A2 _3145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5394__A2 _4318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6591__A1 _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7465__B _2709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7135__A3 _2257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5450_ _0883_ _0887_ _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_121_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6343__A1 as2650.stack\[4\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_25_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9008__CLK clknet_leaf_76_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6894__A2 _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5381_ _0741_ _0772_ _0819_ _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7120_ _2375_ _2385_ _2391_ _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_114_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_2_0_wb_clk_i clknet_0_wb_clk_i clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_141_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8096__A1 _3326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7051_ _2329_ _2332_ _2333_ _1295_ _0163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__6646__A2 _1855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6002_ _1387_ _0717_ _4390_ _1388_ _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_132_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8399__A2 _3582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5004__I _4269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7071__A2 _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7953_ _2338_ _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4843__I _4315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6904_ as2650.r123_2\[1\]\[7\] _2189_ _2203_ _2204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7884_ _3121_ _3123_ _3124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_63_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6835_ _2128_ _2149_ _2150_ _2151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_51_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_64_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6766_ _2082_ _2083_ _2085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4999__B _4370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8505_ _3515_ _3698_ _3701_ _3626_ _3702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5717_ _1140_ _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5674__I _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6697_ _0427_ _1837_ _1819_ _2016_ _2017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_108_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8436_ _0605_ _0619_ _3635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5648_ _1077_ _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5137__A2 _4304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8367_ _1484_ _0458_ _3567_ _3568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_30_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6885__A2 _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5579_ _1012_ _0012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7318_ _2466_ _2576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8087__A1 _3313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8298_ _2712_ _2748_ _3501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_104_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7834__A1 _2869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7249_ _1407_ _2513_ _2514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7834__B2 _2735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output36_I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5073__A1 _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5073__B2 _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8225__I _3435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4820__A1 _4238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8562__A2 _3754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7117__A3 _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6325__A1 _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8078__A1 _3277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7732__C _2758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7825__A1 _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4928__I _4415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4639__A1 _4218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput8 io_in[8] net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_76_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8563__C _2437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8250__A1 _2284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5064__A1 _4193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4950_ _0388_ _0392_ _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_45_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8002__A1 _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4881_ _0323_ _0324_ _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_75_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8553__A2 _3731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6620_ as2650.r0\[6\] _4381_ _1935_ _0466_ _1942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_60_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6564__A1 _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7761__B1 _3004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6551_ _4210_ _4321_ _0832_ _1874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8305__A2 _3503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7108__A3 _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5502_ net10 _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6482_ _1804_ _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8221_ _1794_ _3412_ _3433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5433_ _0870_ _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4878__A1 _4356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8069__A1 _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8152_ _1363_ _3379_ _2586_ _3380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5364_ _0802_ _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7103_ _1343_ _1452_ _1453_ _2374_ _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__6619__A2 _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8083_ as2650.psu\[3\] _3252_ _0936_ _3315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5295_ _0734_ _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7034_ _2316_ _1462_ _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7292__A2 _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7044__A2 _2324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8241__A1 as2650.stack\[7\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8985_ _0146_ clknet_leaf_3_wb_clk_i as2650.r123_2\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5669__I _4289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8792__A2 _3940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7936_ _3172_ _3173_ _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_36_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7867_ _2732_ _3106_ _3107_ _3087_ _3108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_54_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8544__A2 _3739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6818_ _2127_ _2134_ _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_7798_ _3029_ _3031_ _3037_ _3039_ _3040_ _3041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_50_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6749_ _2013_ _2067_ _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6307__A1 _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8419_ _2910_ _3618_ _3492_ _3619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4869__A1 _4178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5530__A2 _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8480__A1 _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5294__A1 _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5294__B2 _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5833__A3 _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7035__A2 _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7586__A3 as2650.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8783__A2 _3940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6794__A1 _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5597__A2 _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5349__A2 _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_35_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6203__I _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8299__A1 _1496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6849__A2 _2151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5521__A2 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4658__I _4238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4875__A4 _4236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5080_ _4012_ _0520_ _0521_ _4002_ _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_97_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7026__A2 _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8223__A1 _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8990__CLK clknet_leaf_68_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6785__A1 _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8770_ _1355_ _3253_ _3939_ _3941_ _3942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_5982_ _4164_ _4099_ _1368_ _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_64_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7982__B1 _3208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7721_ _2775_ _2965_ _1471_ _2966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4933_ _0374_ _0375_ _0371_ _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8526__A2 _3058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7652_ _2897_ _2898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_61_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6537__A1 _1859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4864_ _4337_ _4345_ _4334_ _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_127_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6603_ _1873_ _1902_ _1925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5438__B _4291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7583_ _2829_ _2830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4795_ _4229_ _4375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_59_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_59_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6113__I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6534_ _0864_ _1843_ _1806_ _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5760__A2 _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6465_ as2650.stack\[1\]\[6\] _1769_ _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5416_ _0828_ _0854_ _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8204_ _1721_ _3419_ _3421_ _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6396_ as2650.pc\[6\] _1737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_47_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4571__I0 _4148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8135_ _0873_ _3362_ _3363_ _3364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5347_ _0718_ _0719_ _0679_ _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8462__A1 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8066_ _1173_ _3252_ _0936_ _3299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5278_ _4397_ _0615_ _0583_ _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_60_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7017_ _2303_ _2304_ _2305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7017__A2 _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8214__A1 _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6776__A1 _2071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8968_ _0129_ clknet_leaf_2_wb_clk_i as2650.r123_2\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7919_ _2736_ _3157_ _3158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8899_ _0060_ clknet_3_3_0_wb_clk_i as2650.psl\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6528__A1 _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6023__I _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8659__B _3842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5862__I _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8863__CLK clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5503__A2 _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6700__A1 _2018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6179__B _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8453__A1 _2868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6059__A3 _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5267__A1 _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6693__I _2012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8205__A1 as2650.stack\[7\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8756__A2 _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4490__A2 _4070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7964__B1 _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5990__A2 _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7192__A1 _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4580_ _4160_ _4161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5742__A2 _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6868__I _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7473__B _2469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5772__I _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6250_ _0981_ _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__7495__A2 _2742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8692__A1 _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5201_ _0636_ _0641_ _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6181_ _1542_ _1557_ _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8444__A1 _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5132_ _0571_ _0573_ _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_112_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5063_ _0490_ _0504_ _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8822_ _2506_ _3978_ as2650.psl\[1\] _3988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5012__I _4276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6758__A1 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5025__A4 _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8753_ _1237_ _2676_ _1424_ _3925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5965_ _4037_ _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5947__I _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5430__A1 _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8323__I _3479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7704_ _1281_ _2860_ _2949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4916_ _4252_ _0346_ _0359_ _4203_ _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_8684_ _0713_ _3840_ _3862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5896_ _1280_ _1290_ _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_139_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5981__A2 _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7635_ _1638_ _2880_ _2881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7183__A1 _4301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4847_ _0290_ _4127_ _4130_ _4132_ _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_7566_ _2735_ _2802_ _2812_ _2813_ _2814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4778_ _4161_ _4237_ _4357_ _4358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__8886__CLK clknet_leaf_52_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5733__A2 _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4536__A3 _4116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6517_ _4045_ _4061_ _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7497_ _1550_ _2600_ _2734_ _2745_ _2746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_134_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6448_ _1772_ _1778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_79_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7891__C1 _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9167_ net46 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6379_ _1721_ _1722_ _1723_ _1724_ _0100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_103_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7830__C _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7238__A2 _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8118_ _3345_ _3346_ _3347_ _3282_ _3348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_103_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9098_ _0259_ clknet_leaf_48_wb_clk_i as2650.stack\[4\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8049_ _3247_ _3283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6018__I _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6749__A1 _2013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7410__A2 _2658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5857__I _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5421__A1 _4138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5724__A2 _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_4_wb_clk_i clknet_3_0_0_wb_clk_i clknet_leaf_4_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_67_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5488__A1 _4129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7229__A2 _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4463__A2 _4043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7401__A2 _2651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5767__I _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4671__I _4226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5750_ _1103_ _1163_ _1165_ _0030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5963__A2 _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4701_ _4259_ _4274_ _4279_ _4280_ _4281_ _4282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_5681_ _1109_ _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7165__A1 _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7420_ _2376_ _2669_ _2670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4632_ _4212_ _4213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7915__C _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6912__A1 as2650.r123_2\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5715__A2 _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7180__A4 _4123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7351_ _2605_ _2607_ _2608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4563_ _4026_ _4143_ _4144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6302_ _1664_ _1665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8665__A1 _3836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7282_ _1550_ _4122_ _2541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7468__A2 _2708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4494_ _4064_ _4074_ _4075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9021_ _0182_ clknet_leaf_7_wb_clk_i as2650.holding_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6233_ _1603_ _1604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6140__A2 _4294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8417__A1 _3596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6164_ _1541_ _0068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8417__B2 _3602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4846__I _4125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5115_ _0292_ _0556_ _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6095_ _1214_ _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_44_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7222__I _2489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5100__B1 _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5046_ _4114_ _0425_ _0487_ _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__7640__A2 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8481__C _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8805_ _1506_ _3969_ _3971_ _3973_ _2639_ _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6997_ _4029_ _1054_ _2275_ _4102_ _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
Xclkbuf_leaf_74_wb_clk_i clknet_3_0_0_wb_clk_i clknet_leaf_74_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_8736_ _1311_ _3906_ _3909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5948_ _1334_ _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8667_ _3838_ _2014_ _3848_ _3849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5879_ _1249_ _1266_ _1270_ _1273_ _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_107_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7618_ _2863_ _2810_ _2864_ _2865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6903__A1 _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8598_ net38 net51 _3716_ _3718_ _3791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__9064__CLK clknet_leaf_39_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7549_ _2796_ _2777_ _2797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8105__B1 _2651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7459__A2 _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6667__B1 _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6131__A2 _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8408__A1 _3603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4693__A2 _4272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8901__CLK clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7092__B1 _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5080__C _4002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7395__A1 _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6198__A2 _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7147__A1 _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7698__A2 _2904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_15_wb_clk_i_I clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6370__A2 _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6211__I _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8647__A1 _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6107__C1 _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6122__A2 _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5881__A1 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4666__I _4244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7042__I _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6920_ _0965_ _1799_ _2218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6851_ _2165_ _2166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5497__I _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6189__A2 _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5802_ _1200_ _1197_ _1202_ _0045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_54_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6782_ _0591_ _1909_ _2099_ _2100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8521_ net35 _3717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__9087__CLK clknet_leaf_26_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5733_ _1110_ _1150_ _1154_ _0024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8452_ _3626_ _3629_ _3650_ _3294_ _3651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_104_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5664_ _1093_ _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7403_ _2647_ _2611_ _2653_ _2654_ _2334_ _2655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_117_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4615_ _4193_ _4195_ _4196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8383_ _3500_ _3583_ _3519_ _3584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5595_ as2650.r123\[0\]\[6\] _0878_ _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_102_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6121__I as2650.psl\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4546_ _4126_ _4127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7334_ _2461_ _2591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8757__B _2706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7310__A1 _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4477_ as2650.idx_ctrl\[0\] _4058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_46_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7265_ _0689_ _2526_ _2500_ _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__8924__CLK clknet_leaf_30_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9004_ _0165_ clknet_leaf_23_wb_clk_i net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6216_ _1587_ _0074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7196_ _2260_ _2466_ _2467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5872__A1 _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8048__I _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6147_ _1518_ _1468_ _1533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6078_ _4037_ _1453_ _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_2
XANTENNA__8810__A1 _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5029_ _0414_ _4319_ _4416_ _0332_ _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_113_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xwrapped_as2650_57 io_oeb[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_68 io_oeb[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xwrapped_as2650_79 io_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_53_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5200__I _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8719_ _0640_ _0355_ _3892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7129__A1 as2650.halted vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6888__B1 _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5356__B _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8667__B _3848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7301__A1 _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7852__A2 _3092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8801__A1 _3911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7797__I _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7368__A1 _2623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6206__I _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5918__A2 _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7135__A4 _2343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7540__A1 _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8947__CLK clknet_leaf_34_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7037__I _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5380_ _0744_ _0771_ _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_126_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8096__A2 _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7050_ net24 _2329_ _2333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6001_ _0346_ _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7952_ _3168_ _3177_ _3189_ _2688_ _3190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_83_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6903_ _0857_ _2012_ _2203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7359__A1 _2613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7883_ _3089_ _3122_ _3123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6116__I net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6834_ _2131_ _2132_ _2129_ _2150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_62_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8020__A2 _2700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5909__A2 _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6031__A1 _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6765_ _2082_ _2083_ _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5955__I _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6582__A2 _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8504_ _3596_ _3700_ _3701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7375__C _2326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5716_ as2650.pc\[14\] _1089_ _1097_ as2650.r123_2\[0\]\[6\] _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__4593__A1 as2650.psl\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6696_ _0431_ _1910_ _2015_ _1821_ _2016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_8435_ _3604_ _3632_ _3605_ _3633_ _3634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_104_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5647_ _4297_ _1075_ _1076_ _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_136_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8366_ _3540_ _3541_ _3566_ _3567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5542__B1 _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5578_ _0999_ _1011_ _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_85_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7391__B _2611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7317_ _1549_ _2450_ _2574_ _2575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5690__I _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4529_ _4016_ _4110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8087__A2 _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8297_ _2559_ _3500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9102__CLK clknet_leaf_13_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7834__A2 _3066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7248_ _2280_ _2513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7179_ _2282_ _2449_ _2450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_24_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7598__A1 _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8547__B1 _3738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output29_I net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5865__I _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4584__A1 _4163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7522__A1 _2759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8078__A2 _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6089__A1 _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput9 io_in[9] net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_76_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4944__I as2650.holding_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8250__A2 _2266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5064__A2 _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4880_ _0300_ _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7761__A1 _2996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7761__B2 _2823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4575__A1 _4113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6550_ _1871_ _0853_ _1872_ _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5501_ _0935_ _0936_ _0938_ _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_118_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6481_ _4131_ _1798_ _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8220_ _1648_ _3419_ _3432_ _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5432_ _0869_ _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_69_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4878__A2 _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8069__A2 _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8151_ _1480_ _3378_ _3379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5363_ _0800_ _0801_ _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7102_ _4005_ _1451_ _1217_ _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_47_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5294_ _0454_ _0600_ _0704_ _0512_ _0733_ _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_8082_ _4206_ _3249_ _3314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_141_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5827__A1 _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7033_ _1271_ _1278_ _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5015__I _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7044__A3 _2326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8241__A2 _3436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8984_ _0145_ clknet_leaf_3_wb_clk_i as2650.r123_2\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5055__A2 _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8792__A3 _2488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7935_ _1128_ _1373_ _3173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7866_ _2779_ _3094_ _2996_ _2770_ _3107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_51_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6004__A1 _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6817_ _2130_ _2133_ _2134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7797_ _2536_ _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8061__I _3269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6748_ _1803_ _2065_ _2066_ _2067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7504__A1 _2710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6679_ _1940_ _1955_ _2000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6307__A2 _1662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8418_ _2851_ _3598_ _3618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_87_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8349_ _3549_ _3550_ _4097_ _3551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_3_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7405__I _4131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5118__I0 as2650.r123\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5294__A2 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6491__A1 _4196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8232__A2 _3437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5046__A2 _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7991__A1 _2561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6794__A2 _2076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6546__A2 _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8471__A2 _3644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7251__S _2501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8223__A2 _3419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5981_ _1240_ _1241_ _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6785__A2 _1966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7982__A1 _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7982__B2 _2689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7720_ _2591_ _2963_ _2964_ _2931_ _2965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_80_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4932_ _0371_ _0374_ _0375_ _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_52_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7651_ _2545_ _2897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4863_ _0297_ _0306_ _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__7734__A1 _2843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6537__A2 _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6602_ as2650.r123_2\[2\]\[1\] _1865_ _1924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7582_ _2683_ _2829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4794_ _4373_ _4374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6533_ _4133_ _1799_ _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6464_ _1789_ _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8203_ _1670_ _3415_ _3420_ _3409_ _3421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5415_ _0830_ _0853_ _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__4849__I _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6395_ _1734_ _1722_ _1735_ _1736_ _0104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7225__I _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8134_ _2036_ _0873_ _3363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4720__A1 _4296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5346_ _0784_ _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4571__I1 _4149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8065_ as2650.overflow _3249_ _3298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_130_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5277_ _0716_ _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6473__A1 _1654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7016_ _2293_ _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7670__B1 _2836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5901__C _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5028__A2 _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8967_ _0128_ clknet_leaf_80_wb_clk_i as2650.r123_2\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6776__A2 _2094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7973__A1 _2462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4787__A1 _4024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7918_ _3139_ _3141_ _3157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_93_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8898_ _0059_ clknet_3_4_0_wb_clk_i as2650.psl\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_54_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7849_ _3054_ _3057_ _3090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__7725__A1 as2650.pc\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6528__A2 _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8150__A1 _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6974__I _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8453__A2 _3631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6059__A4 _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5267__A2 _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_62_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7964__A1 _2857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7964__B2 _2882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7738__C _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6214__I _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7192__A2 _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7246__S _2501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4950__A1 _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8141__A1 _3338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8692__A2 _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5200_ _0504_ _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6180_ _1556_ _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5131_ _0572_ _0474_ _0573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6455__A1 _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5258__A2 _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5062_ _4191_ _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_57_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6207__A1 _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8821_ _1777_ _2504_ _3986_ _3987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7955__A1 _2830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6758__A2 _2076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8752_ _2664_ _3923_ _3924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4769__A1 _4326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5964_ _1348_ _1349_ _1350_ _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7007__I0 _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7703_ _4095_ _2416_ _2948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4915_ _0349_ _0354_ _0358_ _4226_ _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_8683_ _3859_ _3836_ _3861_ _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7707__A1 _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5895_ as2650.psu\[5\] _1283_ _1286_ _1289_ _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_61_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7634_ _1684_ _2833_ _2880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_138_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4846_ _4125_ _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7183__A2 _4084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8380__A1 _3537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5194__A1 _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7565_ _2745_ _2813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4777_ _4161_ _4356_ _4276_ _4357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6516_ _1838_ _1839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4941__A1 _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7496_ _1255_ _2708_ _2745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4579__I _4152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6447_ _4377_ _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8683__A2 _3836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9166_ net46 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7891__B1 _3117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6378_ _1615_ _1718_ _1719_ _1724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8495__B _2482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8117_ _0875_ _2960_ _3347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5329_ _0747_ _0761_ _0768_ _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_130_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9097_ _0258_ clknet_leaf_54_wb_clk_i as2650.stack\[4\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8048_ _0934_ _3282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6997__A2 _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8199__A1 _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7246__I0 _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7839__B _2927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6749__A2 _2067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6743__B _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5359__B _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6034__I _4049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6969__I _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5185__A1 _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4932__A1 _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8123__A1 _2431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8674__A2 _3846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8980__CLK clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6685__A1 _2003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5488__A2 _4312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6918__B _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6988__A2 _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4999__A1 _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6653__B _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7937__A1 _2788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7401__A3 _2652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_44_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5412__A2 _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6460__I1 _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5963__A3 _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4700_ _4135_ _4281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5680_ _1106_ _1090_ _1098_ as2650.r123_2\[0\]\[1\] _1108_ _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XANTENNA__8362__A1 net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7165__A2 _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5176__A1 _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4631_ _4001_ as2650.ins_reg\[1\] _4212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_50_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6912__A2 _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7350_ _2550_ _2606_ _2595_ _2607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_15_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4562_ _4069_ _4143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8114__A1 _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6301_ _1663_ _1605_ _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8665__A2 _3845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7281_ _2341_ _2321_ _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4493_ _4025_ as2650.ins_reg\[7\] _4074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5479__A2 _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6676__A1 _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9020_ _0181_ clknet_leaf_8_wb_clk_i as2650.holding_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6232_ _1602_ _1147_ _1603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6828__B _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8417__A2 _3598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6163_ as2650.r123_2\[3\]\[7\] _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6428__A1 _1646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7625__B1 _2849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5114_ _4368_ _0516_ _0555_ _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6428__B2 as2650.stack\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6094_ _1479_ _0782_ _1480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_100_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5100__B2 _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5045_ as2650.holding_reg\[4\] _4114_ _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5651__A2 _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7928__A1 _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8804_ _3869_ _0803_ _3972_ _3973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_20_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6996_ _4091_ _2286_ _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_53_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6600__A1 _4355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8735_ _1311_ _3906_ _3907_ _3908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5947_ _1091_ _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8666_ _1619_ _3843_ _3848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8353__A1 _3472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5878_ _1272_ _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7617_ _0429_ _0340_ _2864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5167__A1 _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4829_ _4370_ _4374_ _4408_ _4409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9165__I net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8597_ _3787_ _3789_ _3472_ _3790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6903__A2 _2012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_43_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_43_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4914__A1 _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7548_ _2444_ _2796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8105__A1 _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8105__B2 _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7479_ _1765_ _2688_ _2728_ _2729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6667__A1 _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6667__B2 _4209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6419__A1 _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6419__B2 as2650.stack\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7092__A1 _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7092__B2 as2650.r123\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7919__A1 _2736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8592__A1 _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7395__A2 _2647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8344__A1 _3540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7147__A2 _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6370__A3 _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6107__B1 _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8647__A2 _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6107__C2 _4242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5108__I _4267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5552__B _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5881__A2 _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7083__A1 _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8876__CLK clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5633__A2 _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_0_wb_clk_i_I clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6850_ _1051_ _1766_ _2165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_78_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8583__A1 _2546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5801_ as2650.stack\[1\]\[9\] _1201_ _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5397__A1 _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6781_ _0602_ _1968_ _1838_ _2098_ _2099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_95_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8520_ net36 _3716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5732_ as2650.stack\[5\]\[9\] _1153_ _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7926__C _2684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8451_ _3537_ _3631_ _3649_ _2580_ _3650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_31_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5663_ _1091_ _1092_ _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7402_ _4048_ _2641_ _2654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6897__A1 as2650.r123_2\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4614_ _4043_ _4194_ _4195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8382_ _2846_ _3582_ _3583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_102_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5594_ _1013_ _0942_ _1026_ _0013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7333_ _1293_ _2590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8638__A2 _3823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4545_ _4064_ _4026_ _4069_ _4126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_102_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6649__A1 _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7264_ _2524_ _2525_ _2526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4476_ as2650.idx_ctrl\[1\] _4057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_144_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7310__A2 _2464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9003_ _0164_ clknet_3_3_0_wb_clk_i net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6215_ _1586_ _1573_ _1557_ _1459_ _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4857__I _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7195_ _2282_ _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7233__I _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5872__A2 _4300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6146_ _1474_ _1476_ _1477_ _1478_ _1531_ _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_97_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7074__A1 _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8810__A2 _3974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6077_ _1463_ _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_3307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6821__A1 _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5028_ _0373_ _0370_ _0470_ _4187_ _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_72_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input10_I wb_rst_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4592__I as2650.carry vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_58 io_oeb[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_69 io_oeb[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7377__A2 _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8574__A1 _2298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5388__A1 _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6979_ _1059_ _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__9031__CLK clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8718_ _0407_ _0412_ _3891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8326__A1 _2803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7129__A2 _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8649_ _1214_ _2319_ _3833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5560__A1 _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5560__B2 _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7301__A2 _2439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5312__A1 _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7143__I _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8899__CLK clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8683__B _3861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7065__A1 _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8565__A1 _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7540__A2 _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5551__A1 as2650.r123\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7481__C _2730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7053__I _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6000_ _0304_ _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input2_I io_in[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8593__B _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7951_ _1008_ _2842_ _3176_ _3187_ _3188_ _3189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_67_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9054__CLK clknet_leaf_64_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6902_ _2147_ _2186_ _2202_ _0145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_36_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7882_ as2650.pc\[9\] _1371_ _3122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8556__A1 _3097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6833_ _2127_ _2134_ _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_62_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6031__A2 _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6764_ _4209_ _0526_ _2083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8308__A1 _4391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8503_ net35 _3699_ _3700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_50_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5715_ _1104_ _1138_ _1139_ _0021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4593__A2 _4173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6695_ _0436_ _1823_ _2015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_13_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6132__I as2650.psl\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8434_ _0539_ _0515_ _3633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5646_ _4003_ _0528_ _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8365_ _0347_ _0321_ _0326_ _3566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__5971__I _4362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5577_ _0558_ _0871_ _0963_ _1010_ _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_7316_ _4036_ _4054_ _2574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4528_ _4108_ _4109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8296_ _1613_ _3491_ _3497_ _3498_ _3499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_105_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5192__B _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7295__A1 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4587__I _4167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7247_ _2512_ _0180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4459_ _4039_ _4040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_137_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7178_ _4036_ _4122_ _2449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7047__A1 _4089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6129_ _4005_ _1514_ _1482_ _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_100_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7598__A2 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8795__A1 _2832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8795__B2 _3920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8547__A1 _3051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5781__A1 _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4584__A2 _4164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7138__I _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6977__I _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6089__A2 _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9077__CLK clknet_leaf_52_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7038__A1 _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8786__A1 _3951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6217__I _4188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5121__I as2650.r0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8538__A1 _3731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8002__A3 _3233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8914__CLK clknet_leaf_33_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4960__I _4299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7761__A2 _2968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4575__A2 _4153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7048__I _2330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5500_ _0937_ _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_125_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6480_ _1802_ _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8710__A1 _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5431_ _0860_ _0868_ _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5791__I _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8150_ _1479_ _1366_ _3377_ _3378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5362_ as2650.holding_reg\[7\] _0716_ _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__8100__C _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7101_ _0462_ _2151_ _2373_ _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_142_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8081_ _3281_ _3313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5293_ _0318_ _0706_ _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_141_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7032_ _1336_ _1223_ _1363_ _1226_ _2315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_99_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5827__A2 _4099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8983_ _0144_ clknet_leaf_3_wb_clk_i as2650.r123_2\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7934_ _3121_ _3169_ _3171_ _3172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8529__A1 _3667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7865_ _0959_ _2961_ _3094_ _3105_ _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__5966__I _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6004__A2 _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8342__I _4060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6816_ _2131_ _2132_ _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7796_ _3038_ _3039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6747_ _0511_ _1832_ _2066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6678_ _1982_ _1998_ _1999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7504__A2 _2749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8701__A1 _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5629_ _4050_ as2650.cycle\[4\] _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8417_ _3596_ _3598_ _3601_ _3602_ _3616_ _3617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_3_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8348_ _1403_ _0331_ _3550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_30_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8465__B1 _3493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5118__I1 as2650.r123_2\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8279_ _2494_ _2571_ _3483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8517__I _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6491__A2 _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output41_I net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5876__I _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5203__B1 _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8153__C1 _2651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5825__B _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7259__A1 _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8456__B1 _3653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8427__I _2580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8759__A1 _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7431__A1 _2401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5980_ _1364_ _0705_ _1366_ _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_65_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7982__A2 _2690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4931_ _0332_ _0373_ _4320_ _0372_ _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XTAP_3490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5993__A1 _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7650_ _1688_ _2880_ _2896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_61_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4862_ _4328_ _0305_ _4344_ _4340_ _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_36_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7734__A2 _2975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6601_ _1905_ _1922_ _1923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_60_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7581_ _2774_ _2828_ _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4793_ _4160_ _4332_ _4372_ _4373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_140_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6532_ _1854_ _1855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7498__A1 _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6463_ _1788_ _1022_ _1778_ _1789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_134_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8202_ as2650.stack\[7\]\[1\] _3412_ _3420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5414_ _0834_ _0836_ _0852_ _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__6410__I _1748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6394_ _1693_ _1717_ _1711_ _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_8133_ _0880_ _3004_ _3361_ _3362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5345_ _0783_ _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4720__A2 _4299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8064_ _3273_ _0316_ _3294_ _3296_ _3297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_99_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5276_ _0715_ _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7015_ _1407_ _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_68_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_68_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6473__A2 _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7670__A1 as2650.stack\[7\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7422__A1 _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8966_ _0127_ clknet_leaf_81_wb_clk_i as2650.r123_2\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7973__A2 _3208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7917_ _1121_ _3155_ _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__4787__A2 _4366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8897_ _0058_ clknet_leaf_50_wb_clk_i as2650.stack\[0\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7848_ _1088_ _1371_ _3089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5736__A1 as2650.stack\[5\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7779_ _2970_ _2974_ _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7489__A1 _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8021__B _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8150__A2 _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6320__I _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7413__A1 _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9115__CLK clknet_leaf_42_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_34_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7964__A2 _3197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_42_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7754__C _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4702__A2 _4186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5130_ _0473_ _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_96_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4685__I as2650.addr_buff\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_73_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6455__A2 _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5061_ _0501_ _0502_ _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_81_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_77_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6207__A2 _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8820_ _1572_ _2504_ _3911_ _3986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7955__A2 _3190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8751_ _2669_ _3923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5963_ _0711_ _0589_ _0517_ _0414_ _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_80_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4769__A2 _4191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8106__B _3276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7007__I1 _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7702_ _2710_ _2947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4914_ _0354_ _0357_ _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8682_ _3838_ _0646_ _3839_ _3860_ _3861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5894_ _1287_ _1288_ _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7707__A2 _2931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7945__B _3182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7633_ _2830_ _2877_ _2879_ _0199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4845_ _4324_ _4412_ _0289_ _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_21_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5718__A1 as2650.r123\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8380__A2 _3564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7564_ _1575_ _2804_ _2808_ _2811_ _2812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4776_ _4057_ as2650.idx_ctrl\[0\] _4356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__6391__A1 _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6515_ _1817_ _1838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7495_ _2594_ _2742_ _2743_ _2606_ _2744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4941__A2 _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7236__I _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6446_ _1614_ as2650.stack\[1\]\[1\] _1769_ _1776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6143__A1 _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8776__B _2534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9165_ net46 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7891__A1 _3039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7891__B2 _3029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6377_ as2650.stack\[3\]\[1\] _1715_ _1723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8116_ as2650.psl\[5\] _3248_ _0886_ _3346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5328_ _0667_ _0767_ _0768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9096_ _0257_ clknet_leaf_53_wb_clk_i as2650.stack\[4\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_138_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8047_ _1267_ _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5259_ _0299_ _0698_ _0486_ _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_87_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6997__A3 _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7246__I1 _2511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7946__A2 _3155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8949_ _0110_ clknet_leaf_34_wb_clk_i as2650.stack\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5709__A1 _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5185__A2 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6382__A1 _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5375__B _4164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8123__A2 _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7331__B1 _2535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5488__A3 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4696__A1 _4275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7634__A1 _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6988__A3 _2266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7749__C _2869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7937__A2 _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6225__I as2650.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5963__A4 _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8362__A2 net53 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8440__I _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4630_ _4210_ _4022_ _4211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5176__A2 _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6373__A1 _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4561_ _4141_ _4142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__7056__I _4284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8114__A2 _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6300_ _0910_ _1296_ _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7280_ _4292_ _2538_ _2539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_144_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4492_ _4063_ _4073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6231_ _1601_ _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6162_ _1540_ _0067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7625__A1 _2647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5113_ _4367_ _0549_ _0554_ _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_69_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7625__B2 _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6093_ _4072_ _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4439__A1 _4018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5044_ _4325_ _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5100__A2 _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5651__A3 _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8803_ _1475_ _3906_ _3972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_93_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6995_ _4047_ _4051_ _2270_ _2271_ _2286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_81_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8734_ _0692_ _0701_ _3907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5946_ as2650.psl\[1\] _0803_ _1328_ _4396_ _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_59_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8665_ _3836_ _3845_ _3847_ _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5877_ _1271_ _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8353__A2 _3554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7616_ _1402_ _4384_ _2863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4828_ _4377_ _4201_ _4369_ _4407_ _4408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5167__A2 _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8596_ _3143_ _2482_ _3788_ _3789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_7547_ _1622_ _2794_ _2795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4914__A2 _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4759_ _4162_ _4169_ _4339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8105__A2 _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7478_ _2438_ _2726_ _2727_ _2728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7864__A1 _3039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6429_ _1642_ _1758_ _1762_ _0112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_136_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4678__A1 _4189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_12_wb_clk_i clknet_3_2_0_wb_clk_i clknet_leaf_12_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_134_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7616__A1 _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9079_ _0240_ clknet_leaf_65_wb_clk_i as2650.stack\[7\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7092__A2 _2054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7919__A2 _3157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8041__A1 _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8041__B2 _3275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8592__A2 _3144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7395__A3 _2611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4602__A1 _4168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5884__I _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8260__I _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6107__A1 _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8647__A3 _2411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6929__B _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7855__A1 _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6658__A2 _1978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7604__I _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4669__A1 _4248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5330__A2 _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7607__A1 _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5881__A3 _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7083__A2 _4315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6830__A2 _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4841__A1 _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8032__A1 _3244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8583__A2 _3770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5800_ _1195_ _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6780_ _1281_ _1910_ _2097_ _1836_ _2098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_90_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6594__A1 _4230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7495__B _2743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5731_ _1148_ _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_95_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5794__I _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8450_ _3638_ _3648_ _3579_ _3649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5662_ _4129_ _0529_ _0884_ _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__8103__C _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7401_ _4261_ _2651_ _2652_ _2653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4613_ _4075_ _4194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8381_ _1621_ _1402_ _3534_ _3582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6897__A2 _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5593_ _0946_ _1024_ _1025_ _1026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_15_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7332_ _1252_ _2589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8099__A1 _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4544_ _4124_ _4125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6649__A2 _1837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7263_ _1584_ _2513_ _2525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4475_ _4055_ _4056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_89_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9002_ _0163_ clknet_leaf_15_wb_clk_i net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6214_ _1393_ _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7194_ _2464_ _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6145_ _1480_ _1530_ _1396_ _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8271__A1 _2606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6076_ _4101_ _1418_ _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8810__A3 _3975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4873__I _4367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5027_ _0467_ _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_59 io_oeb[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8970__CLK clknet_leaf_34_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5388__A2 _4321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6978_ _4051_ _2269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8717_ _0639_ _2096_ _3890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5929_ _0501_ _0627_ _1315_ _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_110_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8326__A2 _3527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7129__A3 _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8648_ _0940_ _2571_ _2673_ _3832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__6337__A1 _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8579_ _3088_ _3740_ _3773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4899__A1 _4218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5560__A2 _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7837__A1 _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7837__B2 _3077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5312__A2 _4415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8262__A1 _3465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8255__I _3458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8565__A2 _3484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6576__A1 _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5119__I _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5303__A2 _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8253__A1 _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5067__A1 _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8993__CLK clknet_leaf_69_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7950_ _2760_ _3168_ _3188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4814__A1 _4064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8005__A1 _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6901_ _0774_ _1905_ _2193_ as2650.r123_2\[1\]\[6\] _2202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_78_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8005__B2 _2656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7881_ _3090_ _3088_ _3121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6832_ _2013_ _2135_ _2147_ _1852_ _2148_ _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_91_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6763_ _0710_ _2036_ _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7509__I _2724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8502_ net34 net52 _3630_ _3699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_108_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6413__I _1751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5714_ as2650.stack\[3\]\[13\] _1086_ _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6694_ _4390_ _2014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8433_ _0538_ _0515_ _3632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5645_ as2650.ins_reg\[3\] _4067_ _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8364_ _3465_ _3565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5576_ _1000_ _0966_ _0930_ _1009_ _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5542__A2 _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7315_ _2263_ _2539_ _2573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4868__I _4168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4527_ _4083_ _4108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8295_ _2472_ _3498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8492__A1 _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7246_ _0387_ _2511_ _2501_ _2512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4458_ as2650.ins_reg\[3\] _4039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7177_ _1568_ _2446_ _2447_ _2418_ _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_8_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8244__A1 _2675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7047__A2 _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6128_ _1508_ _1510_ _1513_ _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_105_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5699__I _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8795__A2 _3962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6059_ _1442_ _1263_ _1278_ _1445_ _1446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XTAP_3127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4805__A1 _4212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8547__A2 _3558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5230__A1 _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5081__I1 as2650.r123_2\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5781__A2 _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7863__B _2433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8866__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5297__A1 _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7038__A2 _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5049__A1 _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7103__B _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6797__A1 _4210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6942__B _2237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5221__A1 _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6233__I _1603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7265__S _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5430_ _0861_ _0867_ _4134_ _4117_ _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__8710__A2 _2522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6721__A1 _4208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5361_ _0799_ _4222_ _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_114_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7100_ _0817_ _2362_ _2368_ as2650.r123\[2\]\[7\] _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8474__A1 _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8080_ _3268_ _0413_ _3270_ _3311_ _3312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_82_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5292_ _4370_ _0709_ _0731_ _0317_ _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_99_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5288__A1 _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7031_ _1272_ _1421_ _2314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9021__CLK clknet_leaf_7_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6408__I _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8982_ _0143_ clknet_leaf_81_wb_clk_i as2650.r123_2\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6788__A1 _2096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4638__I1 as2650.r123\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_fanout53_I net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7933_ _3089_ _3122_ _3148_ _3170_ _3171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__7948__B _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5460__A1 _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7864_ _3039_ _3096_ _3104_ _2465_ _3105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_110_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6815_ _2120_ _2118_ _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6004__A3 _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7795_ _2548_ _2466_ _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7239__I _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6746_ _0516_ _2056_ _2064_ _2065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8889__CLK clknet_leaf_64_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5763__A2 _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6960__A1 _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6677_ _1985_ _1997_ _1998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_109_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8701__A2 _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8416_ _3609_ _3615_ _3515_ _3616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5628_ _4120_ _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_136_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8347_ _3510_ _3511_ _3548_ _3549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_133_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5559_ _0987_ _0990_ _0993_ _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_69_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8465__A1 _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7268__A2 _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8278_ _3462_ _3474_ _3481_ _1473_ _3482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8465__B2 _3662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7229_ _1797_ _1436_ _1440_ _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7702__I _2710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8217__A1 _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6318__I _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6779__A1 _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7976__B1 _3211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_24_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output34_I net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5451__A1 _4290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_3_1_0_wb_clk_i clknet_0_wb_clk_i clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5203__A1 _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6053__I _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5203__B2 _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6951__A1 _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5754__A2 _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5892__I _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8153__C2 _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5825__C _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9044__CLK clknet_leaf_29_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8456__A1 _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7259__A2 _2521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8456__B2 _3654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6937__B _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8759__A2 _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6228__I _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7431__A2 _2452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4971__I _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4930_ _0333_ _4320_ _0372_ _0373_ _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_80_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5993__A2 _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4861_ _4326_ _0304_ _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6600_ _4355_ _1803_ _1921_ _1922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_61_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5745__A2 _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4792_ _4160_ _4371_ _4269_ _4372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7580_ _2775_ _2827_ _1471_ _2828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6531_ _1853_ _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8695__A1 _2307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6462_ _1645_ as2650.stack\[1\]\[5\] _1767_ _1788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_140_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8201_ _3409_ _3419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5413_ _0841_ _0851_ _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_127_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6393_ as2650.stack\[3\]\[5\] _1731_ _1735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5344_ net3 _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8132_ _1492_ _3248_ _3360_ _0879_ _3361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_126_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4720__A3 _4300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4571__I3 _4151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8063_ _2623_ _0331_ _3295_ _2547_ _3296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5275_ _4211_ _4216_ _4220_ _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_87_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7014_ _2293_ _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7422__A2 _2325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8965_ _0126_ clknet_leaf_76_wb_clk_i as2650.r123_2\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5977__I _4224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7916_ _3111_ _3083_ _3067_ _3155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
Xclkbuf_leaf_37_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_102_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8896_ _0057_ clknet_leaf_51_wb_clk_i as2650.stack\[0\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7186__A1 _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7847_ _3082_ _2987_ _3088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5736__A2 _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6933__A1 _1978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7778_ _1650_ _1373_ _3021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9067__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6729_ _1987_ _2048_ _2049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_20_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7489__A2 _2703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8150__A3 _3377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_30_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7860__C _3100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7110__A1 _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7661__A2 _2858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5672__A1 _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5672__B2 as2650.r123_2\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8610__A1 net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5887__I _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5424__A1 _4111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6621__B1 _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7177__A1 _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6924__A1 _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8429__A1 _2933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7101__A1 _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7342__I _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5060_ _0388_ _0383_ _0392_ _0497_ _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_112_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5663__A1 _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7404__A2 _4048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8750_ _1228_ _1250_ _2335_ _3922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_19_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5962_ _0333_ _4376_ _4188_ _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_20_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7701_ _1287_ _2868_ _2869_ _2945_ _2946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4913_ _0355_ _0356_ _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_8681_ _0590_ _3840_ _3860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5893_ _4310_ _1245_ _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_90_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7632_ _1729_ _2878_ _2339_ _2879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7945__C _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4844_ as2650.r123\[1\]\[1\] _4413_ _0287_ _0288_ _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6915__A1 _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7563_ _2809_ _2810_ _2811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_105_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6391__A2 _1712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4775_ _4354_ _4355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_105_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6514_ _1836_ _1837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7494_ _1400_ _2416_ _2743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7961__B _2708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6445_ _1775_ _0115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7340__A1 _2449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8927__CLK clknet_leaf_39_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_9164_ net46 net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7891__A2 _3115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6376_ _1711_ _1722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8115_ as2650.psu\[5\] _3251_ _3345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5327_ _0762_ _0763_ _0766_ _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_87_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9095_ _0256_ clknet_leaf_55_wb_clk_i as2650.stack\[4\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8140__I0 _3368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7643__A2 _2848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8046_ _3268_ _4355_ _3270_ _3279_ _3280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_88_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5258_ _0689_ _0680_ _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5189_ _0495_ _0498_ _0629_ _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8948_ _0109_ clknet_leaf_34_wb_clk_i as2650.stack\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_73_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8879_ _0040_ clknet_leaf_58_wb_clk_i as2650.stack\[2\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_12_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6906__A1 _1842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5709__A2 _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7331__A1 _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7331__B2 _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4696__A2 _4276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5893__A1 _4310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7162__I _2433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7634__A2 _2833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8831__A1 _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6988__A4 _2278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7398__A1 _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6070__A1 _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8362__A3 net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7337__I _2593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7570__A1 as2650.stack\[7\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6241__I _1610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4560_ _4140_ _4141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4491_ _4063_ _4068_ _4071_ _4072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_143_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6230_ _0861_ _1600_ _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_87_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8168__I _3389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6161_ as2650.r123_2\[3\]\[6\] _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5112_ _4264_ _0553_ _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7625__A2 _2834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6092_ _1362_ _1397_ _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5636__A1 _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4439__A2 _4019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5043_ _4324_ _0461_ _0485_ _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8802_ _1474_ _3970_ _3969_ _3971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6994_ _4105_ _1845_ _2285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8733_ as2650.holding_reg\[7\] _2493_ _3905_ _3906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5945_ _1329_ _1331_ _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8664_ net42 _3846_ _3847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_107_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5876_ _1069_ _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7615_ _2861_ _2862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4827_ _4378_ _4406_ _4407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8595_ _3144_ _3728_ _3788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7546_ _1613_ _2703_ _2794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4758_ _4156_ _4157_ _4338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_120_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7477_ _2683_ _2727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4689_ _4267_ _4269_ _4270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_107_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9105__CLK clknet_leaf_13_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6428_ _1646_ _1759_ _1760_ as2650.stack\[2\]\[5\] _1755_ _1762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_134_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7864__A2 _3096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5875__A1 _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6359_ _1707_ _0097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7616__A2 _4384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8813__A1 _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9078_ _0239_ clknet_leaf_51_wb_clk_i as2650.stack\[7\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_52_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_52_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_8029_ _1464_ _3264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_76_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_17_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8041__A2 _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8592__A3 _3765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7866__B _2996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8329__B1 _3530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7552__A1 _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7304__A1 _4194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6107__A2 _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4669__A2 _4249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7607__A2 _2834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8804__A1 _3869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4841__A2 _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6236__I _1606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7791__A1 _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7495__C _2606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5730_ _1103_ _1150_ _1152_ _0023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_128_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5661_ _4083_ _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8740__B1 _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7400_ _4128_ _2273_ _2652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_90_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4612_ _4192_ _4193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8380_ _3537_ _3564_ _3580_ _2629_ _3581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_117_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5592_ _0651_ _0870_ _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7331_ _1551_ _2572_ _2588_ _2535_ _2275_ _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_116_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4543_ _4118_ _4123_ _4124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7262_ _1028_ _1286_ _2524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4474_ _4050_ as2650.cycle\[4\] _4052_ _4054_ _4055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
X_9001_ _0162_ clknet_leaf_12_wb_clk_i as2650.addr_buff\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6213_ _1585_ _0073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_132_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7193_ _1546_ _2464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6144_ _1383_ _1366_ _1529_ _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_86_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8271__A2 _2469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6075_ _4260_ _4108_ _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6282__A1 _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5026_ _0468_ _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4832__A2 _4355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5050__I _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6977_ _1450_ _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7782__A1 _2843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8361__I net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4596__A1 as2650.psl\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8716_ _3595_ _3889_ _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5928_ _0800_ _0801_ _0682_ _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8647_ _2253_ _2317_ _2411_ _3831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_5859_ _4032_ _1253_ _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_107_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8578_ _3763_ _3768_ _3771_ _2629_ _3772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_108_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4899__A2 _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7529_ _1622_ _2776_ _2777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7837__A2 _2961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4520__A1 _4070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8262__A2 _4279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7440__I _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7470__B1 _2719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6056__I _4105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6576__A2 _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7525__A1 _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7615__I _2861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5839__A1 as2650.psl\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4974__I _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5067__A2 _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4814__A2 _4248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6900_ _2107_ _2192_ _2201_ _0144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_48_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7880_ _3119_ _3120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_63_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6831_ as2650.r123_2\[2\]\[6\] _2069_ _2148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7764__A1 _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6762_ _2079_ _2080_ _2081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_62_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8501_ _3691_ _3692_ _3696_ _3697_ _3698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_50_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5713_ _1137_ _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6693_ _2012_ _2013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8432_ net52 _3630_ _3631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5644_ _1073_ _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8363_ _3562_ _3563_ _3564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5575_ _0966_ _1008_ _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7314_ _2571_ _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4526_ _4086_ _4098_ _4106_ _4107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__4750__A1 _4325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8294_ _3496_ _3497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_117_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7245_ _2509_ _2510_ _2511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4457_ _4037_ _4038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8492__A2 _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7176_ _1251_ _0888_ _1094_ _1465_ _2447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_28_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6127_ _1511_ _4392_ _0539_ _4015_ _1512_ _1513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__8244__A2 _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6058_ _1251_ _1444_ _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_46_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_14_wb_clk_i_I clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4805__A2 _4384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5009_ _0451_ _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_73_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6007__A1 _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7507__A1 _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5518__B1 _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8180__A1 _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8040__B _3270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7435__I _2684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_53_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6494__A1 _4202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8235__A2 _3440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7443__B1 _2692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7994__A1 _4133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6797__A2 _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5221__A2 _4318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4980__A1 _4218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6721__A2 _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4732__A1 _4311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5360_ as2650.holding_reg\[7\] _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_127_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8474__A2 _3572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5291_ _0713_ _4201_ _4258_ _0730_ _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__8960__CLK clknet_leaf_43_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5288__A2 _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7030_ _2313_ _0162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8981_ _0142_ clknet_leaf_0_wb_clk_i as2650.r123_2\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7985__A1 _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7932_ _1120_ _1491_ _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5460__A2 _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7863_ _3101_ _3103_ _2433_ _3104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7737__A1 _2979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6814_ _2113_ _2117_ _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6424__I _1748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7794_ _2558_ _2594_ _3034_ _3036_ _3037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5212__A2 _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6745_ _1808_ _2062_ _2063_ _2064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_56_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6676_ _1989_ _1996_ _1997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_109_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8162__A1 _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8415_ _1411_ _3509_ _3614_ _2626_ _3615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5627_ _4118_ _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8346_ _1502_ _4374_ _3548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5558_ as2650.stack\[6\]\[11\] _0952_ _0992_ _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4509_ _4046_ _4090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8277_ _2473_ _3478_ _3480_ _1667_ _3481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8465__A2 _2975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5489_ _4313_ _0926_ _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5279__A2 _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7228_ _1358_ _1551_ _1562_ _2496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_120_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7159_ _2430_ _2431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7976__A1 _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7976__B2 _3029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5451__A2 _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output27_I net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7728__A1 _2933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6400__A1 _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8153__A1 _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8983__CLK clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8456__A2 _3480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_7_wb_clk_i clknet_3_2_0_wb_clk_i clknet_leaf_7_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_2_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6509__I _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7967__A1 _2462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7431__A3 _2618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6244__I _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5288__C _4204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4860_ _4332_ _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_2791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8392__A1 _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8392__B2 _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4791_ _4268_ as2650.addr_buff\[5\] _4371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6530_ _1822_ _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8144__A1 _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4699__I _4273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6461_ _1787_ _0119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8695__A2 _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7498__A3 _2734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8200_ _1709_ _3410_ _3414_ _3418_ _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5412_ _0847_ _0850_ _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_115_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6392_ _0590_ _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8131_ _1375_ _3248_ _3360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_142_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5343_ _4206_ _4379_ _4174_ _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_138_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6458__A1 as2650.stack\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8062_ _2256_ _0327_ _3295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5274_ _0537_ _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7013_ as2650.addr_buff\[3\] _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_114_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7958__A1 _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8964_ _0125_ clknet_leaf_76_wb_clk_i as2650.r123_2\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6630__A1 _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8856__CLK clknet_leaf_55_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7915_ _2947_ _3150_ _3153_ _1285_ _3154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_36_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8895_ _0056_ clknet_leaf_51_wb_clk_i as2650.stack\[0\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7846_ _3084_ _3086_ _3087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7186__A2 _2456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_77_wb_clk_i clknet_3_0_0_wb_clk_i clknet_leaf_77_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_75_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7777_ as2650.pc\[7\] net2 _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_71_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4989_ _4226_ _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7591__C1 _2836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6728_ _2034_ _2047_ _2048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_137_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8135__A1 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8686__A2 _3839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6659_ as2650.r123_2\[2\]\[2\] _1865_ _1980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__9117__D _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6697__A1 _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8329_ _1622_ _3525_ _3530_ _2473_ _3531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_105_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7949__A1 _2813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6621__A1 _4382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7177__A2 _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8374__A1 _3549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6924__A2 _2213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8677__A2 _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7101__A2 _2151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5112__A1 _4264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8879__CLK clknet_leaf_58_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6860__A1 _1611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5663__A2 _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4982__I _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4915__C _4226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6612__A1 _4376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5415__A2 _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6463__I1 _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5961_ _4294_ _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_98_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_3_2_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7700_ _2942_ _2944_ _2945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_59_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4912_ _4395_ _4398_ _4238_ _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_8680_ net19 _3859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_34_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5892_ _1281_ _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8365__A1 _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7631_ _2683_ _2878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5179__A1 _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4843_ _4315_ _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6915__A2 _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7562_ _2805_ _2807_ _2810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_105_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8117__A1 _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4774_ _4330_ _4353_ _4354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_144_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8122__C _2724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6513_ _1820_ _1836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8668__A2 _3846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7493_ _2740_ _2741_ _2742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_140_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7961__C _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6444_ _1771_ _4306_ _1774_ _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7340__A2 _2596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8629__I _3819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6375_ _1610_ _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8114_ _1365_ _0591_ _3344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5326_ as2650.r0\[0\] _0765_ _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9094_ _0255_ clknet_leaf_51_wb_clk_i as2650.stack\[4\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8140__I1 _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8045_ _3277_ _4374_ _3278_ _3273_ _3279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5103__A1 _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5257_ _4172_ _0685_ _0696_ _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5053__I _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7689__B _2933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5188_ _0628_ _0493_ _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4862__B1 _4344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4892__I _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8364__I _3465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6603__A1 _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8947_ _0108_ clknet_leaf_34_wb_clk_i as2650.stack\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__9034__CLK clknet_leaf_41_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8356__A1 _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8878_ _0039_ clknet_leaf_58_wb_clk_i as2650.stack\[2\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_40_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7829_ _2321_ _3071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8313__B _3515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6906__A2 _1911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8659__A2 _3836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5590__A1 _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7331__A2 _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5893__A2 _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7095__A1 _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5898__I _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7398__A2 _2650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8595__A1 _3144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6070__A2 _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6522__I _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4908__A1 _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5581__A1 as2650.stack\[3\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4490_ _4026_ _4070_ _4071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6160_ _1539_ _0066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5111_ _0552_ _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7086__A1 _4283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6091_ _1340_ _1346_ _1356_ _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_112_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8822__A2 _3978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5636__A2 _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5042_ as2650.r123\[1\]\[3\] _4304_ _0484_ _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9057__CLK clknet_leaf_66_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7389__A2 _2637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8801_ _3911_ _2510_ _2509_ _3970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6993_ _1567_ _2282_ _1430_ _2283_ _2284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_19_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6061__A2 _1447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5944_ as2650.psl\[1\] _0803_ _1330_ _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8732_ _2493_ _1340_ _3905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8663_ _3835_ _3846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5875_ _1269_ _1222_ _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7614_ _2860_ _2861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4826_ _4379_ _4380_ _4405_ _4406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8594_ _3785_ _3786_ _3506_ _3787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7545_ _0883_ _2736_ _2793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4757_ _4334_ _4336_ _4337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5048__I as2650.holding_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7476_ _1667_ _2689_ _2690_ _2700_ _2725_ _2726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4688_ _4268_ as2650.addr_buff\[5\] _4269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8510__A1 _3702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6427_ _1636_ _1758_ _1761_ _0111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_108_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5875__A2 _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6358_ as2650.r123\[3\]\[6\] _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_1_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7077__A1 net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5309_ _0664_ _0747_ _0748_ _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_9077_ _0238_ clknet_leaf_52_wb_clk_i as2650.stack\[7\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6289_ _1040_ _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8813__A2 _3975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5088__B1 _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6824__A1 _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8028_ _1462_ _3263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5511__I _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8577__A1 _3505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4555__C _4135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6052__A2 _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8592__A4 _3766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7866__C _2770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8329__A1 _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8329__B2 _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7438__I _2687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7001__A1 _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6342__I _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7552__A2 _2787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8501__A1 _3691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7304__A2 _4056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_opt_2_0_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4797__I _4376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7068__A1 _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8568__A1 _3595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8032__A3 _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8917__CLK clknet_leaf_33_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7240__A1 _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_23_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7791__A2 _2991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5577__B _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6252__I as2650.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5660_ _1089_ _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__8740__A1 _3303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4611_ _4191_ _4192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_129_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5591_ _0966_ _1021_ _1023_ _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_106_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7330_ _1569_ _2578_ _2583_ _2480_ _2587_ _2588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_102_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4542_ _4119_ _4122_ _4123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_117_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7261_ _2523_ _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4473_ _4053_ _4033_ _4054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_132_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9000_ _0161_ clknet_leaf_10_wb_clk_i as2650.addr_buff\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6212_ _1584_ _1576_ _1557_ _1243_ _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_125_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7192_ _1459_ _1460_ _2456_ _2463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_135_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7059__A1 _4166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6143_ _1481_ _1525_ _1526_ _1528_ _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6074_ _1242_ _1459_ _1460_ _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7032__B _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5025_ _4375_ _4187_ _0370_ _0467_ _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_6_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7967__B _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6976_ _1421_ _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_54_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7782__A2 _3024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8715_ as2650.psl\[5\] _3882_ _3888_ _3889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5927_ _0511_ _0650_ _1313_ _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__4596__A2 as2650.carry vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5858_ _1061_ _1246_ _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_8646_ net41 _3830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_16_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4809_ _4388_ _4389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__4979__S0 _4002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8577_ _3505_ _3770_ _3771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_5789_ _0890_ _0897_ _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7528_ _1612_ _1597_ _2776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7298__A1 _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7459_ _4243_ _2415_ _2285_ as2650.addr_buff\[0\] _2709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_108_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_43_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5950__B _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8798__A1 _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5156__S0 _4003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7470__A1 _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5241__I _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7470__B2 _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5481__B1 _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_60_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7168__I _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6072__I _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8722__A1 _4325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5839__A2 _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4898__I0 as2650.r123\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7631__I _2683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7461__A1 as2650.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5151__I as2650.r0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7213__A1 _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6830_ _1964_ _2146_ _2147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6761_ _2041_ _2043_ _2080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8500_ _1393_ _3565_ _3464_ _3697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5712_ _1135_ _1090_ _1098_ as2650.r123_2\[0\]\[5\] _1136_ _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_56_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6692_ _1963_ _2012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8713__A1 _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8431_ net32 _3597_ _3630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5643_ _4063_ _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8362_ net30 net53 net28 _3563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5574_ _1004_ _1007_ _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8130__C _3269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7313_ _2277_ _2571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4525_ _4039_ _4101_ _4105_ _4106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_8293_ _3040_ _2749_ _3493_ _3495_ _3496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_85_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7244_ _2299_ _1286_ _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4456_ _4031_ _4036_ _4037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7175_ _2445_ _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_67_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7541__I _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6126_ _1375_ _0725_ _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7452__A1 _1597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6057_ _4361_ _1443_ _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_46_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5463__B1 _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5008_ _0443_ _0400_ _0446_ _0447_ _0450_ _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_73_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5996__I _4072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6007__A2 _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7204__A1 _2336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7204__B2 _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5766__A1 _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6959_ _2162_ _2207_ _2227_ _2250_ _2251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_126_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5010__B _4273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8704__A1 _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7507__A2 _2755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5518__A1 as2650.stack\[2\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8629_ _3819_ _3820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8321__B _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7716__I _2823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8180__A2 _3398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7691__A1 _2891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6494__A2 _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7451__I _2469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7443__A1 as2650.stack\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7443__B2 as2650.stack\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__9118__CLK clknet_leaf_46_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7994__A2 _2676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6797__A3 _2042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5757__A1 _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_3_7_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5855__B _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4980__A2 _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5347__S _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4732__A2 _4312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5146__I _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5290_ _4378_ _0729_ _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4985__I _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7682__A1 _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8980_ _0141_ clknet_leaf_2_wb_clk_i as2650.r123_2\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7931_ _3119_ _3147_ _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4638__I3 as2650.r123_2\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7862_ _2793_ _3102_ _3103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7737__A2 _2980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6813_ _2128_ _2129_ _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7793_ _2897_ _3035_ _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7964__C _3200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6744_ _0553_ _1966_ _2063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6675_ _1991_ _1995_ _1996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_91_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8162__A2 _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5626_ _4102_ _1055_ _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8414_ _3509_ _3613_ _3614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7980__B _3208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8345_ _1404_ _3544_ _3507_ _3547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5557_ _0915_ _0991_ _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4508_ _4088_ _4089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8276_ _3479_ _3480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5488_ _4129_ _4312_ _0529_ _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7673__A1 _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5279__A3 _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7227_ _1214_ _0397_ _1345_ _2495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4439_ _4018_ _4019_ _4020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7271__I _2530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7158_ _1242_ _2430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7425__A1 _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6109_ _0400_ _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8622__B1 _3813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7089_ _4317_ _2010_ _2364_ as2650.r123\[2\]\[2\] _2367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7976__A2 _2979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5739__A1 _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6400__A2 _1712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8138__C1 _3264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8153__A2 _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7664__A1 _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7967__A2 _2782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__9090__CLK clknet_leaf_24_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7431__A4 _2680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4790_ _4369_ _4370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8144__A2 _1475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6260__I _1627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6460_ _1786_ _1000_ _1778_ _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5411_ _0844_ _0848_ _0849_ _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_12_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6391_ _1636_ _1712_ _1733_ _0103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8130_ _3324_ _0700_ _3357_ _3358_ _3269_ _3359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_5342_ _0780_ _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_126_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8061_ _3269_ _3294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7655__A1 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5273_ _0712_ _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7012_ _2300_ _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_29_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7407__A1 _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8963_ _0124_ clknet_leaf_77_wb_clk_i as2650.r123_2\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5969__A1 _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7914_ _2796_ _3142_ _3151_ _3152_ _3153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_102_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6630__A2 _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5479__C _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8894_ _0055_ clknet_leaf_52_wb_clk_i as2650.stack\[0\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7845_ _3083_ _3085_ _3086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8383__A2 _3583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5197__A2 _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6394__A1 _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7776_ _3015_ _3018_ _3019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4988_ _0430_ _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7591__B1 _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6727_ _2046_ _2047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_71_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8135__A2 _3362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6170__I _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6146__A1 _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6658_ _1964_ _1978_ _1979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7894__A1 _2470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_46_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_46_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5609_ _1039_ _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6697__A2 _1837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6589_ _4106_ _1805_ _1911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8328_ _2884_ _2787_ _3475_ _3529_ _3530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_117_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8259_ _2405_ _3463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8071__A1 _3303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8046__B _3270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6621__A2 _1935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_62_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8950__CLK clknet_leaf_34_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5188__A2 _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5112__A2 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8062__A1 _2256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6612__A2 _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6255__I _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5960_ _1340_ _0778_ _1346_ _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_46_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4911_ _0324_ _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_94_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5891_ _1285_ _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7630_ _2831_ _2874_ _2876_ _2877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4842_ _0286_ _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5179__A2 _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7561_ _2320_ _2809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4773_ _4331_ _4334_ _4351_ _4352_ _4353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_144_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8117__A2 _2960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6512_ _1801_ _1834_ _1835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6128__A1 _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7492_ _1502_ _4233_ _2741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_101_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6443_ _1773_ _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6374_ _1709_ _1712_ _1716_ _1720_ _0099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_66_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5351__A2 _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8113_ _3341_ _3342_ _3269_ _3343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_103_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5325_ _0764_ _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9093_ _0254_ clknet_leaf_25_wb_clk_i net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_88_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8044_ _3277_ _4359_ _3278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5256_ _4343_ _0688_ _0692_ _0312_ _0695_ _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__6300__A1 _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5187_ _0488_ _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_99_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6593__C _1842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4862__A1 _4328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8053__A1 _4417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6165__I _4006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7800__A1 _2781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6603__A2 _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8973__CLK clknet_leaf_35_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8946_ _0107_ clknet_leaf_33_wb_clk_i as2650.stack\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4614__A1 _4043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8877_ _0038_ clknet_leaf_58_wb_clk_i as2650.stack\[2\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8356__A2 _2490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7828_ _3067_ _3069_ _3070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6367__A1 _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7564__B1 _2808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4917__A2 _4239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7759_ as2650.stack\[2\]\[6\] _1047_ _3000_ _3002_ _3003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_127_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5590__A2 _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7867__A1 _2732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7867__B2 _3087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7331__A3 _2588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7619__A1 _2863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8292__A1 _2804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7095__A2 _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8044__A1 _3277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8595__A2 _3728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4605__A1 _4147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6070__A3 _4202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5030__A1 _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5581__A2 _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7858__A1 _2743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8846__CLK clknet_leaf_69_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5110_ _0550_ _0513_ _0514_ _0447_ _0551_ _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7086__A2 _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6090_ _4127_ _1475_ _1337_ _1476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_111_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5041_ _0462_ _0483_ _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8996__CLK clknet_leaf_23_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4844__A1 as2650.r123\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4844__B2 _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_0_wb_clk_i wb_clk_i clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_8800_ _3873_ _3877_ _3968_ _3969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_93_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6597__A1 _4374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6992_ _4035_ _1062_ _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8731_ _3890_ _3902_ _3903_ _3904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_81_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5943_ _0698_ _0692_ _0802_ _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_34_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8662_ _3838_ _3258_ _3844_ _3845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5874_ _1267_ _1268_ _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7613_ _1072_ _2860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4825_ _4240_ _4404_ _4405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8593_ _3144_ _3766_ _2301_ _3786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7544_ _2780_ _2790_ _2791_ _2792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_33_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4756_ as2650.holding_reg\[1\] _4332_ _4336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4687_ as2650.addr_buff\[6\] _4268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7475_ _2701_ _2721_ _2722_ _2723_ _2724_ _2725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_88_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6426_ _1639_ _1759_ _1760_ as2650.stack\[2\]\[4\] _1755_ _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA_clkbuf_leaf_33_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6521__A1 _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6357_ _1706_ _0096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7077__A2 _2357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8274__A1 _2701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5308_ _0666_ _0667_ _0670_ _0671_ _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__8274__B2 _3477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9076_ _0237_ clknet_leaf_53_wb_clk_i as2650.stack\[7\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6288_ _1649_ _1637_ _1652_ _0081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5999__I _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5088__B2 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8027_ _4379_ _3262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5239_ _0594_ _0596_ _0598_ _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_102_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8026__A1 _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8577__A2 _3770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5013__B _4356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8929_ _0090_ clknet_leaf_32_wb_clk_i as2650.stack\[4\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5260__A1 _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8329__A2 _3525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7001__A2 _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_61_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_61_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_130_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6760__A1 _2037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8869__CLK clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8265__A1 _3468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7068__A2 _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8285__I _3459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4826__A1 _4379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5149__I _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5003__A1 _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8740__A2 _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4610_ _4190_ _4191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5590_ _1022_ _0947_ _0929_ _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5554__A2 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4541_ _4120_ _4121_ _4028_ _4122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__4988__I _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7364__I _2559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4472_ as2650.cycle\[1\] _4053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7260_ _0636_ _2522_ _2500_ _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6503__A1 _4243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9024__CLK clknet_leaf_7_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6211_ _1412_ _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7191_ _2461_ _2462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_125_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6142_ _1527_ _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6073_ _4100_ _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5024_ _0466_ _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7032__C _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5490__A1 _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7231__A2 _2496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6975_ _1443_ _4123_ _2265_ _2266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_81_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6443__I _1773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8714_ _3869_ _3886_ _3882_ _3887_ _3888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5926_ _0700_ _1312_ _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5793__A2 _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8645_ _1211_ _3821_ _3829_ _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5857_ _1251_ _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_55_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4808_ _4383_ _4385_ _4387_ _4388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_4
X_8576_ net38 _3769_ _3770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_107_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5788_ _1102_ _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7527_ _2684_ _2775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4739_ _4319_ _4320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8495__A1 _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7458_ _1079_ _2708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6409_ _1747_ _1177_ _1601_ _1748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_7389_ _2408_ _2637_ _2642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_118_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8247__A1 _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8798__A2 _2677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9059_ _0220_ clknet_leaf_40_wb_clk_i as2650.stack\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_44_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5156__S1 _4013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4808__A1 _4383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7470__A2 _2707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5784__A2 _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8722__A2 _4159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9047__CLK clknet_leaf_30_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8486__A1 _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4898__I1 as2650.r123\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__9051__D _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5432__I _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7997__B1 _1843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7461__A2 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7213__A2 _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8410__A1 _2899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6263__I _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6760_ _2037_ _2042_ _2079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_63_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5711_ _1013_ _4290_ _1094_ _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6691_ _1962_ _1979_ _1980_ _2011_ _0125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__8713__A2 _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8430_ _2932_ _3628_ _3629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5642_ _4124_ _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8361_ net31 _3562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_129_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5573_ _0916_ _1005_ _1006_ _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4511__I _4091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7312_ _1550_ _2535_ _2557_ _2570_ _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_144_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4524_ _4104_ _4105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8292_ _2804_ _3494_ _2750_ _3495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7243_ _0981_ _1348_ _2509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4455_ _4032_ _4035_ _4036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7174_ _2444_ _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8139__B _3359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6125_ as2650.psl\[1\] _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_140_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5342__I _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7978__B _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6056_ _4105_ _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7452__A2 _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8653__I _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5007_ _0448_ _0449_ _4371_ _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7204__A2 _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6173__I _4035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6963__A1 _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6958_ as2650.r123_2\[0\]\[7\] _2223_ _2250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_81_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5909_ as2650.stack\[0\]\[8\] _1302_ _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6889_ _1923_ _2192_ _2194_ _0140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8704__A2 _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8628_ _3818_ _3819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6715__A1 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5518__A2 _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7218__B _2484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8559_ net51 _3753_ _3754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_108_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7691__A2 _2935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7443__A2 _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7994__A3 _2276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5206__A1 _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6954__A1 _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5757__A2 _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6706__A1 _2013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5855__C _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4568__I0 as2650.r123\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8459__A1 net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8738__I _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7131__A1 _4090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5162__I net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7930_ _1129_ _3167_ _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_49_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7861_ _1106_ _3067_ _3102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_36_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6812_ _1986_ _2084_ _2129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_58_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7792_ _3032_ _2991_ _3033_ _3035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__6945__A1 _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6743_ _1000_ _1908_ _1810_ _2061_ _2062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_108_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8698__A1 _2658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6674_ _1993_ _1994_ _1995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_52_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8413_ _1409_ _0553_ _3612_ _3613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__8162__A3 _1750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5625_ _4029_ _1054_ _4119_ _4033_ _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_118_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8344_ _3540_ _3543_ _3545_ _3546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5556_ as2650.stack\[7\]\[11\] _0891_ _0903_ as2650.stack\[4\]\[11\] as2650.stack\[5\]\[11\]
+ _0907_ _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__5920__A2 _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4507_ _4087_ _4088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7122__A1 _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8275_ _1553_ _1547_ _2471_ _3479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_2_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5487_ _0901_ _0917_ _0919_ _0924_ _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_7226_ _1462_ _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_116_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4438_ as2650.ins_reg\[1\] _4019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5684__A1 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7157_ net54 _2428_ _1459_ _2429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_113_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7425__A2 _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8622__A1 _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6108_ _1486_ _1489_ _1493_ _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_101_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8622__B2 _3654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7088_ _4412_ _2361_ _2366_ _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6039_ _4260_ _4291_ _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_58_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5800__I _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7189__A1 _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5739__A2 _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6936__A1 _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8332__B _2786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8138__B1 _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8138__C2 _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8051__C _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7361__A1 _2615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7890__C _3129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6787__B _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7113__A1 _2347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7664__A2 _2809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5427__A1 _4093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4650__A2 as2650.ins_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6927__A1 _1922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7637__I _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7352__A1 _2336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5410_ _0563_ _0524_ _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6390_ as2650.stack\[3\]\[4\] _1731_ _1732_ _1711_ _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_115_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5341_ _4222_ _0443_ _0777_ _0550_ _0779_ _0447_ _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7104__A1 _4049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7655__A2 _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8060_ _1721_ _3276_ _3280_ _3293_ _2639_ _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5272_ _0711_ _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_130_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7011_ _2298_ _2299_ _2294_ _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_99_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8604__A1 _2892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7407__A2 _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6716__I _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8080__A2 _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8962_ _0123_ clknet_leaf_77_wb_clk_i as2650.r123_2\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5969__A2 _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6091__A1 _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_fanout51_I net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7913_ _0431_ _2593_ _2354_ _3152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_37_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8893_ _0054_ clknet_leaf_53_wb_clk_i as2650.stack\[0\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_24_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7844_ _1088_ _3052_ _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8152__B _2586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7775_ _0922_ _3016_ _3017_ _3018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4987_ _0429_ _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6394__A2 _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7591__A1 as2650.stack\[7\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6726_ _2035_ _2045_ _2046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_71_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6657_ _1965_ _1976_ _1977_ _1978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6146__A2 _1476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5608_ _0792_ _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7894__A2 _3131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6588_ _1853_ _1910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8327_ _1405_ _2261_ _3528_ _3529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_121_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5539_ _0968_ _0970_ _0974_ _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_69_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8258_ _2620_ _2713_ _3462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7209_ _2455_ _2477_ _2478_ _2479_ _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__5016__B _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_15_wb_clk_i clknet_3_3_0_wb_clk_i clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_59_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8189_ _1174_ _1298_ _1591_ _3408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_59_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5409__A1 as2650.r0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8071__A2 _3258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output32_I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5896__A1 _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8288__I _3479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8834__A1 _2519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4765__B _4162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7141__B _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8062__A2 _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5820__A1 _4314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8751__I _2669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4910_ _4024_ _0353_ _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5890_ _1284_ _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_94_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4841_ _0284_ _0285_ _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__7367__I _2622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7573__A1 _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7560_ _2805_ _2807_ _2808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4772_ _4141_ _4336_ _4164_ _4352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_140_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6511_ _4186_ _1803_ _1833_ _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7325__A1 _2344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7491_ _4241_ _4151_ _2740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6442_ _1772_ _1773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_23_wb_clk_i_I clknet_opt_3_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8198__I _3408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6373_ _1599_ _1718_ _1719_ _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
Xclkbuf_3_0_0_wb_clk_i clknet_0_wb_clk_i clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_8112_ _2623_ _0587_ _2547_ _3342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7089__B1 _2364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5324_ as2650.r123\[0\]\[6\] as2650.r123_2\[0\]\[6\] as2650.psl\[4\] _0764_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__8825__A1 _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9092_ _0253_ clknet_leaf_26_wb_clk_i net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_114_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8043_ _2622_ _3277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5255_ _0410_ _0694_ _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6874__C _2165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5186_ _0626_ _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4862__A2 _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8053__A2 _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7800__A2 _3011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8945_ _0106_ clknet_leaf_56_wb_clk_i as2650.stack\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_3_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4614__A2 _4194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8876_ _0037_ clknet_leaf_49_wb_clk_i as2650.stack\[2\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_7827_ _3051_ _3068_ _3069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7277__I _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7564__A1 _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6367__A2 _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_62_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6906__A4 _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7758_ _3001_ _3002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_138_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6709_ _2003_ _2005_ _2029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_123_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6119__A2 _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7689_ _2887_ _2889_ _2933_ _2934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8513__B1 _3709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6130__B _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7619__A2 _2810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8816__A1 _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8292__A2 _3494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8044__A2 _4359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7896__B _2770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4605__A2 _4159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7307__A1 _4056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7858__A2 _3098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5869__A1 _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9054__D _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8807__A1 _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6467__S _1778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8283__A2 _3460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6294__A1 as2650.stack\[5\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5040_ _0481_ _0482_ _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4844__A2 _4413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6991_ _2281_ _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7794__A1 _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6597__A2 _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8730_ _0692_ _0701_ _3903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5942_ _1324_ _1316_ _1327_ _1328_ _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_111_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8661_ _1610_ _3843_ _3844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7546__A1 _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5873_ _4073_ _4077_ _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_94_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4514__I as2650.addr_buff\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7612_ _1631_ _2858_ _2859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4824_ _4252_ _4390_ _4403_ _4404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8592_ _2301_ _3144_ _3765_ _3766_ _3785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_7543_ _2460_ _2791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4755_ _4178_ _4298_ _4335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_88_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7474_ _2430_ _2724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4686_ as2650.addr_buff\[6\] _4266_ _4267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6425_ _1751_ _1760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5345__I _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6521__A2 _1843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4532__A1 _4062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6356_ as2650.r123\[3\]\[5\] _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5307_ _0666_ _0667_ _0670_ _0671_ _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8274__A2 _2713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9075_ _0236_ clknet_leaf_54_wb_clk_i as2650.stack\[7\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_62_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8940__CLK clknet_leaf_42_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6287_ _1651_ _1625_ _1616_ as2650.stack\[5\]\[6\] _1593_ _1652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_142_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8026_ _1422_ _3257_ _3260_ _3261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5238_ _4138_ _0651_ _0678_ _0005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6176__I _4105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5169_ _0432_ _0602_ _0609_ _4204_ _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6037__A1 _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8605__B _3151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7785__A1 _2576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4599__A1 _4177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8928_ _0089_ clknet_leaf_32_wb_clk_i as2650.stack\[4\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_71_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5260__A2 _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8859_ _0020_ clknet_leaf_48_wb_clk_i as2650.stack\[3\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4424__I _4004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7001__A3 _2284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_32_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6760__A2 _2042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_30_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_30_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6512__A2 _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8265__A2 _4272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7403__C _2334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6028__A1 _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5251__A2 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7528__A1 _1612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8250__B _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6751__A2 _2069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4540_ as2650.cycle\[2\] _4121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_106_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4762__A1 _4335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4471_ _4051_ _4030_ _4052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8963__CLK clknet_leaf_77_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6210_ _1582_ _1583_ _0072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7190_ _2460_ _2461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6141_ _4078_ _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6267__A1 _1629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6072_ _1344_ _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4817__A2 _4396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5023_ _0465_ _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5490__A2 _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7767__A1 as2650.pc\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6974_ _1079_ _2265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7231__A3 _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4672__C _4252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8144__C _3294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5242__A2 _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5925_ _4186_ _4355_ _0316_ _0412_ _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_8713_ _2481_ _0511_ _3887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7519__A1 _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6990__A2 _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8644_ as2650.stack\[4\]\[14\] _3819_ _3829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5856_ as2650.halted _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8192__A1 _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4807_ _4217_ _4386_ _4387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8575_ net51 net36 _3718_ _3769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_124_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7555__I _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5787_ _1143_ _1181_ _1189_ _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_72_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7526_ _1679_ _2731_ _2774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4753__A1 as2650.holding_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4738_ _4318_ _4319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7457_ _2539_ _2706_ _2707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__8495__A2 _3572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5075__I _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4669_ _4248_ _4249_ _4250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_107_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4505__A1 _4045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6408_ _1173_ _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7388_ _2408_ _2637_ _2641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7504__B _2752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8247__A2 _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6339_ _1651_ _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_66_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5803__I _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6258__A1 _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9058_ _0219_ clknet_leaf_39_wb_clk_i as2650.stack\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_76_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8009_ _3243_ _3244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4419__I net54 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5481__A2 _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6430__A1 _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6430__B2 as2650.stack\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7893__C _2335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8183__A1 _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6733__A2 _2052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8986__CLK clknet_leaf_69_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6497__A1 _4225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8238__A2 _3438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6249__A1 _1611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7446__B1 _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7997__A1 _2860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7997__B2 _4096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5869__B _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7749__A1 _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7213__A3 _2482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8410__A2 _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6421__A1 _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6421__B2 as2650.stack\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5710_ as2650.pc\[13\] _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6690_ _1867_ _2010_ _2011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_31_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5641_ _1069_ _1070_ _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7921__A1 _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8360_ _3338_ _3561_ _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5572_ as2650.stack\[7\]\[12\] _0892_ _0899_ as2650.stack\[6\]\[12\] _1006_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_117_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7311_ _2534_ _2352_ _2568_ _2569_ _2570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_4523_ _4102_ _4030_ _4103_ _4104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_8291_ net53 _3447_ _3494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__8477__A2 _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6488__A1 _4310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7242_ _2503_ _2507_ _2508_ _0179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4454_ _4034_ _4035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7173_ _1224_ _2353_ _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__8229__A2 _3437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5623__I as2650.cycle\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8139__C _3367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6124_ _4173_ _4241_ _0430_ _4207_ _1509_ _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_115_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7988__A1 _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6055_ _1075_ _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_26_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6660__A1 _1941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5463__A2 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8859__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5006_ _0323_ _0324_ _0399_ _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_113_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8155__B _3382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6412__A1 _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6957_ _2246_ _2247_ _2249_ _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_78_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6963__A2 _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5908_ _1300_ _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6888_ _0287_ _1905_ _2193_ as2650.r123_2\[1\]\[1\] _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__8165__A1 _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8627_ _0967_ _1145_ _3818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5839_ as2650.psl\[7\] _0528_ _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7912__A1 _3143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8558_ _3716_ _3718_ _3753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7509_ _2724_ _2758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_135_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8489_ _3489_ _3685_ _3686_ _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8468__A2 _3661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6479__A1 _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7140__A2 _2411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7979__A1 _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8640__A2 _3823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6100__B1 _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6651__A1 _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7994__A4 _3228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6403__A1 _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5206__A2 _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9014__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6954__A2 _2213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4965__A1 _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8156__A1 _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7409__B _2658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7195__I _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4612__I _4192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4568__I1 as2650.r123_2\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5390__A1 _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5142__A1 _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6983__B _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7798__C _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8631__A2 _3821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6642__A1 _4294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7860_ _2947_ _3092_ _3087_ _2599_ _3100_ _3101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_36_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6811_ _1986_ _2082_ _2128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7791_ _3032_ _2991_ _3033_ _3034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_36_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6742_ _1971_ _2060_ _2061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6673_ _0593_ _1951_ _1994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5618__I _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8698__A2 _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5624_ _1053_ _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8412_ _3610_ _3611_ _3612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4708__A1 _4286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8343_ _3540_ _3543_ _3544_ _3545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5555_ as2650.stack\[2\]\[11\] _0920_ _0988_ as2650.stack\[0\]\[11\] _0989_ _0990_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_118_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4506_ _4067_ _4087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8274_ _2701_ _2713_ _3475_ _3477_ _3478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_69_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5486_ as2650.stack\[7\]\[8\] _0893_ _0920_ as2650.stack\[6\]\[8\] _0923_ _0924_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__7122__A2 _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7225_ _0640_ _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_4437_ _4001_ _4018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5353__I _4210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6881__A1 _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5684__A2 _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7156_ _2427_ _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_8_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6107_ _1490_ _0540_ _1491_ _1492_ _0895_ _4242_ _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8622__A2 _3480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7087_ _4317_ _1960_ _2364_ as2650.r123\[2\]\[1\] _2366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6038_ _1421_ _1424_ _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_73_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9037__CLK clknet_leaf_30_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7189__A2 _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7989_ _1243_ _1352_ _2656_ _3224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4947__A1 _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8138__A1 _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7229__B _1440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8689__A2 _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4432__I _4012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5372__A1 _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8310__A1 _3468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5124__B2 _4229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5675__A2 _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6872__A1 _1646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7899__B _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6872__B2 as2650.stack\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8074__B1 _3263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5427__A2 _4091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6624__A1 as2650.r0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7411__C _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8377__A1 _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6927__A2 _2208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4938__A1 _4324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8129__A1 _3340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4770__C _4298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9057__D _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_13_wb_clk_i_I clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5363__A1 _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7653__I _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5340_ _0715_ _0778_ _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_115_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7104__A2 _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8301__A1 _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5115__A1 _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6269__I _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5271_ _0710_ _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7010_ _1405_ _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6863__A1 _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8604__A2 _3150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7407__A3 _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8417__C _3616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5418__A2 _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6615__A1 _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8961_ _0122_ clknet_leaf_56_wb_clk_i as2650.stack\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_49_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6091__A2 _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7912_ _3143_ _2803_ _3151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8892_ _0053_ clknet_leaf_52_wb_clk_i as2650.stack\[0\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_110_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7843_ as2650.pc\[9\] as2650.pc\[8\] _3052_ _3084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_110_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_58_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7040__A1 _4035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_52_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4986_ net8 _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_75_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7774_ as2650.stack\[4\]\[7\] _2819_ _2956_ as2650.stack\[5\]\[7\] _3017_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_51_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7049__B _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6725_ _2040_ _2044_ _2045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6656_ _0316_ _1965_ _1977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8540__A1 _3340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5607_ as2650.r123\[0\]\[7\] _0963_ _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5354__A1 _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6587_ _1818_ _1909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8326_ _2803_ _3527_ _3528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_121_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5538_ as2650.stack\[0\]\[10\] _0971_ _0973_ as2650.stack\[1\]\[10\] _0974_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5106__A1 _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8257_ _2571_ _3461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5469_ _0906_ _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7208_ _1294_ _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8188_ _1698_ _3386_ _3407_ _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_82_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7139_ _0785_ _2409_ _2410_ _2411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_120_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7004__S _2294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5409__A2 _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6606__A1 _1878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_55_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_55_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_98_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6082__A2 _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8359__A1 net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output25_I net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7031__A1 _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8531__A1 _4097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_124_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5207__B _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6845__A1 _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7422__B _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8598__A1 net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5820__A2 _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7648__I _2687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7022__A1 _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4840_ _4377_ _4322_ _4417_ _4189_ _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8770__A1 _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5584__A1 _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4771_ _4342_ _4347_ _4348_ _4350_ _4351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_105_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6510_ _4279_ _1808_ _1831_ _1832_ _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_105_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7490_ _1481_ _2737_ _2738_ _2739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_144_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5336__A1 _4138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6441_ _1146_ _1177_ _1591_ _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__4800__I _4203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6372_ _1710_ _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8111_ _3340_ _0619_ _3341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7089__A1 _4317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5323_ as2650.r0\[2\] _0560_ _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9091_ _0252_ clknet_leaf_25_wb_clk_i net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8825__A2 _4311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6836__A1 _4225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8042_ _3243_ _3276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5254_ _0689_ _0397_ _0403_ _0693_ _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_142_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5185_ _0623_ _0624_ _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_111_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8589__A1 _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8147__C _3282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8589__B2 _3461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7051__C _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8944_ _0105_ clknet_leaf_56_wb_clk_i as2650.stack\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5811__A2 _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8875_ _0036_ clknet_leaf_46_wb_clk_i as2650.stack\[6\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_64_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7826_ _1656_ _3030_ _3068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7564__A2 _2804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6367__A3 _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8761__A1 _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7757_ as2650.stack\[0\]\[6\] _2819_ _2694_ as2650.stack\[1\]\[6\] _3001_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4969_ _4147_ _0384_ _0409_ _0411_ _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_6708_ _2000_ _2001_ _1999_ _2028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_123_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7316__A2 _4054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8513__A1 _1656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7688_ as2650.pc\[4\] net9 _2933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8513__B2 _3654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5327__A1 _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6639_ _1867_ _1960_ _1961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5806__I _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4710__I _4037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8277__B1 _3480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8309_ _3510_ _3511_ _3512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7619__A3 _2864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6827__A1 _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8057__C _2603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5802__A2 _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5030__A3 _4319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8504__A1 _3596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7307__A2 _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5318__A1 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5869__A2 _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4541__A2 _4121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8807__A2 _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8248__B _3451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7491__A1 _4241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7243__A1 _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6990_ _1074_ _1077_ _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7794__A2 _2594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8892__CLK clknet_leaf_52_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5941_ _0800_ _0811_ _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_0_wb_clk_i clknet_3_0_0_wb_clk_i clknet_leaf_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_8660_ _3837_ _3843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5872_ _1073_ _4300_ _4071_ _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__7546__A2 _2703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8743__A1 _3880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7611_ _1621_ _1612_ _2703_ _2858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4823_ _4227_ _4402_ _4403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5557__A1 _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8591_ _3625_ _3783_ _3784_ _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8711__B _3313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7542_ _2782_ _2777_ _2787_ _2788_ _2789_ _2790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
X_4754_ _4333_ _4334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_105_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7473_ _1666_ _1354_ _2469_ _2723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4685_ as2650.addr_buff\[5\] _4266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4780__A2 _4359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7046__C _2254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6424_ _1748_ _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6521__A3 _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6355_ _1705_ _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6885__C _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5306_ _0661_ _0662_ _0745_ _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_9074_ _0235_ clknet_leaf_51_wb_clk_i as2650.stack\[7\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6286_ _1650_ _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5237_ as2650.r123\[1\]\[5\] _4413_ _0677_ _4316_ _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_8025_ _1383_ _3258_ _4224_ _1528_ _3259_ _3260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_130_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5168_ _0605_ _0354_ _0608_ _4227_ _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_124_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6037__A2 _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5099_ _4042_ _4126_ _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8927_ _0088_ clknet_leaf_39_wb_clk_i as2650.stack\[4\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7288__I _2546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6192__I _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4705__I _4014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8858_ _0019_ clknet_leaf_58_wb_clk_i as2650.stack\[3\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7809_ _3050_ _3051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5548__A1 _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8789_ _3950_ _3958_ _3959_ _3659_ _0275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XPHY_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5536__I _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5980__B _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5720__A1 as2650.stack\[3\]\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_70_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_70_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__8068__B _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5271__I _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8515__C _3711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4834__I0 as2650.r123\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7198__I _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7528__A2 _1597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4470_ as2650.cycle\[6\] _4051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6140_ _0792_ _4294_ _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7464__A1 _2710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6277__I as2650.pc\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6071_ _4109_ _4225_ _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5181__I _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5022_ _0464_ _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7216__A1 _4095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7767__A2 as2650.pc\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6973_ _4044_ _1052_ _2263_ _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__9070__CLK clknet_leaf_41_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8712_ _3313_ _0681_ _3885_ _3886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5924_ _0804_ _0815_ _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_94_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8716__A1 _3595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7519__A2 _2767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8643_ _1209_ _3821_ _3828_ _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_61_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5855_ _1232_ _1245_ _1227_ _1249_ _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_61_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8192__A2 _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4806_ as2650.r123\[1\]\[2\] as2650.r123\[0\]\[2\] as2650.r123_2\[1\]\[2\] as2650.r123_2\[0\]\[2\]
+ _4018_ _4011_ _4386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_8574_ _2298_ _3767_ _3768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5786_ as2650.stack\[2\]\[14\] _1179_ _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7525_ _2640_ _2773_ _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_120_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4737_ _4149_ _4318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4753__A2 _4332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7456_ _1254_ _2282_ _2706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4668_ _4161_ _4249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4505__A2 _4061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6407_ _1745_ _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7571__I _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7387_ _2639_ _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4599_ _4177_ _4158_ _4179_ _4180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7504__C _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6338_ as2650.stack\[4\]\[6\] _1677_ _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5091__I as2650.r0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9057_ _0218_ clknet_leaf_66_wb_clk_i as2650.r0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6269_ _1635_ _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8008_ _3242_ _3243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7207__A1 net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_44_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8707__A1 _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6981__A3 _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8183__A2 _3398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6650__I _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5941__A1 _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7694__A1 _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4898__I3 as2650.r123_2\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7446__B2 as2650.stack\[5\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7997__A2 _4396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8526__B _3721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9093__CLK clknet_leaf_25_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4680__A1 _4260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7749__A2 _2868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7213__A4 _2325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7656__I _2901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5640_ _4170_ _4044_ _4214_ _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5571_ as2650.stack\[4\]\[12\] _0988_ _0972_ as2650.stack\[5\]\[12\] _1005_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_129_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5932__A1 _4159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4522_ as2650.cycle\[1\] as2650.cycle\[0\] _4103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_129_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7310_ _1560_ _2464_ _2569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8290_ _3492_ _3493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6488__A2 _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4453_ _4033_ _4034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_105_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7241_ _4326_ _2503_ _2508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5696__B1 _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7172_ net49 _2426_ _2443_ _1295_ _0174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_125_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6123_ as2650.psl\[7\] _1499_ _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6054_ _4007_ _1440_ _1245_ _1441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_39_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7340__B _2434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5005_ _4265_ _0304_ _4388_ _0344_ _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_22_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8155__C _2730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6412__A2 _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6956_ _2146_ _2229_ _2227_ _2248_ _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_82_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5907_ _1300_ _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6887_ _2188_ _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_70_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8626_ _3625_ _3816_ _3817_ _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5838_ as2650.psl\[6\] _4004_ _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7912__A2 _2803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8557_ _3464_ _3749_ _3751_ _2256_ _3752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__5923__A1 _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5086__I _4019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5769_ _1174_ _1177_ _1084_ _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_120_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7508_ _2744_ _2746_ _2747_ _2756_ _2757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_136_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8488_ net34 _3523_ _3191_ _3686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6479__A2 _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7676__A1 as2650.stack\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7439_ _1423_ _2689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7007__S _2294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5687__B1 _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7428__A1 _2676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9109_ _0270_ clknet_leaf_9_wb_clk_i as2650.ins_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6100__A1 _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7600__A1 _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8953__CLK clknet_leaf_59_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6403__A2 _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4965__A2 _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8156__A2 _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7903__A2 _3141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7667__A1 _2909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7131__A3 _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5142__A2 _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7419__A1 _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8616__B1 _3807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6890__A2 _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6983__C _4284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8092__A1 _3277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7160__B _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6642__A2 _4301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4653__A1 _4212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6810_ _2111_ _2123_ _2126_ _2127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_42_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7790_ net3 _4215_ _3033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_51_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6741_ _1388_ _1909_ _2059_ _2060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8147__A2 _3019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6290__I _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6672_ _1990_ _1992_ _1993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_52_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8698__A3 _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8411_ _2899_ _0451_ _3549_ _3573_ _3574_ _3611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_5623_ as2650.cycle\[2\] _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_104_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4708__A2 _4288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8342_ _4060_ _3544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5554_ as2650.stack\[1\]\[11\] _0972_ _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7658__A1 _2900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4505_ _4045_ _4061_ _4085_ _4086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_8273_ _3447_ _2546_ _3476_ _3477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5485_ _0922_ _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4678__C _4258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8010__I _3244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4436_ _4015_ _4016_ _4017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7224_ _2488_ _2491_ _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5133__A2 _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7155_ _0883_ _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8083__A1 as2650.psu\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6106_ net27 _1492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_140_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7086_ _4283_ _2361_ _2365_ _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_81_wb_clk_i_I clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7830__A1 _3063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8976__CLK clknet_leaf_58_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6037_ _1255_ _1422_ _1223_ _1423_ _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__7830__B2 _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4644__A1 _4080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7988_ _2331_ _3221_ _3222_ _3223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6939_ _0994_ _2213_ _2221_ _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5809__I _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8138__A2 _3263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4713__I _4293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8609_ _3796_ _3801_ _3485_ _3802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5372__A2 _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4869__B _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7649__A1 _2882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8310__A2 _3512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6321__A1 _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8074__A1 _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8074__B2 _2014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8076__B _3308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6375__I _1610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4635__A1 _4214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8377__A2 _3572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4938__A2 _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8129__A2 _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5060__A1 _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4623__I _4203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7888__A1 _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8849__CLK clknet_leaf_67_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5454__I _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8301__A2 _3465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5270_ _0593_ _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_9_wb_clk_i_I clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6312__A1 _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8765__I _2603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6285__I as2650.pc\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8960_ _0121_ clknet_leaf_43_wb_clk_i as2650.stack\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7911_ _3147_ _3149_ _3150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_55_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8891_ _0052_ clknet_leaf_51_wb_clk_i as2650.stack\[0\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8714__B _3882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8368__A2 _3568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7842_ _3082_ _3083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_58_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6379__A1 _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7040__A2 _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7773_ as2650.stack\[7\]\[7\] _2762_ _1046_ as2650.stack\[6\]\[7\] _3016_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4985_ _0427_ _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5051__A1 _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4533__I _4113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6724_ _2041_ _2043_ _2044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_137_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6655_ _0327_ _1907_ _1975_ _1976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5606_ _1037_ _0014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6551__A1 _4210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6586_ _1842_ _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8325_ net30 _3526_ _3527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_106_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5537_ _0972_ _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8256_ _3459_ _3460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5468_ _0905_ _0897_ _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_87_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9004__CLK clknet_leaf_23_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7207_ net25 _2455_ _2478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4419_ net54 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_8_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8187_ _1741_ _3388_ _3390_ as2650.stack\[6\]\[7\] _3384_ _3407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_114_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5399_ as2650.r0\[5\] _0367_ _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_115_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8056__A1 _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7138_ _2394_ _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7803__A1 _2779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7069_ _1226_ _2349_ _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4617__A1 _4196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8359__A2 _3460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7031__A2 _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5042__A1 as2650.r123\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output18_I net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_24_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_24_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4599__B _4179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5274__I _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7098__A2 _2364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6845__A2 _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4856__A1 _4383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4618__I _4198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5281__A1 _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5820__A3 _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7022__A2 _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5033__A1 _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5449__I _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7573__A3 _2820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6781__A1 _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4770_ _4192_ _4239_ _4349_ _4298_ _4350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6440_ _1765_ _1768_ _1770_ _1771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5336__A2 _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6533__A1 _4133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9027__CLK clknet_leaf_17_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6371_ _1717_ _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8110_ _2626_ _3340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7089__A2 _2010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5322_ as2650.r0\[1\] _0523_ _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9090_ _0251_ clknet_leaf_24_wb_clk_i net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8825__A3 _3975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8041_ _1709_ _3245_ _3267_ _3275_ _2590_ _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__6836__A2 _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5253_ _0397_ _0601_ _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4847__A1 _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5184_ _0623_ _0624_ _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6229__B _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4528__I _4108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8943_ _0104_ clknet_leaf_37_wb_clk_i as2650.stack\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_95_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8874_ _0035_ clknet_leaf_46_wb_clk_i as2650.stack\[6\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8210__A1 as2650.stack\[7\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7825_ _1088_ _1655_ _3030_ _3067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_52_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8761__A2 _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7756_ _0949_ _2999_ _3000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_40_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6772__A1 _2028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5575__A2 _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4968_ _0410_ _0382_ _4146_ _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6707_ as2650.r123_2\[2\]\[3\] _1865_ _2027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7687_ as2650.pc\[5\] net1 _2932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_2
X_4899_ _4218_ _0342_ _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6638_ _1927_ _1930_ _1959_ _1960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__6524__A1 _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6569_ _4382_ _0526_ _0845_ _4375_ _1892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5094__I _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8277__A1 _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8308_ _4391_ _4373_ _3511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8277__B2 _1667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8239_ as2650.stack\[7\]\[13\] _3436_ _3445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5822__I _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4838__A1 _4376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4438__I as2650.ins_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5263__A1 _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5269__I _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6212__B1 _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6763__A1 _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5030__A4 _4416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4901__I _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7712__B1 _2956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4829__A1 _4370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8248__C _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7491__A2 _4151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7243__A2 _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4792__B _4269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5940_ _1315_ _1326_ _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_93_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5871_ _1265_ _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5006__A1 _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7610_ _2704_ _2857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4822_ _4393_ _4245_ _4401_ _4402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8590_ net38 _3713_ _3714_ _3784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6754__A1 _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7541_ _1273_ _2789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4753_ as2650.holding_reg\[1\] _4332_ _4333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_109_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5907__I _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4811__I net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7472_ _2427_ _2713_ _2722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4684_ _4153_ _4265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6423_ _1745_ _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6354_ as2650.r123\[3\]\[4\] _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8439__B _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5305_ _0418_ _0372_ _0565_ _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_9073_ _0234_ clknet_leaf_38_wb_clk_i as2650.stack\[7\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5642__I _4124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6285_ as2650.pc\[6\] _1650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8024_ _2349_ _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5236_ _0676_ _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5493__A1 _4306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5493__B2 _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5167_ _0354_ _0607_ _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8431__A1 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6037__A3 _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5098_ _0539_ _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_44_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7785__A3 _3027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8926_ _0087_ clknet_leaf_32_wb_clk_i as2650.stack\[4\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6993__A1 _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8857_ _0018_ clknet_leaf_57_wb_clk_i as2650.stack\[3\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__8734__A2 _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7808_ as2650.pc\[8\] _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8788_ _0902_ _3950_ _3959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7739_ _2576_ _2978_ _2982_ _2983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_36_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8498__A1 _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4771__A3 _4348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7170__A1 _2438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4523__A3 _4103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8349__B _4097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5720__A2 _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7473__A2 _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8422__A1 _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5501__B _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6383__I _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5787__A2 _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4834__I1 as2650.r123_2\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6736__A1 _1962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5727__I _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_opt_3_1_wb_clk_i_I clknet_opt_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5711__A2 _4290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7464__A2 _2713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8661__A1 _1610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6070_ _1343_ _1091_ _4202_ _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5475__A1 _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_input9_I io_in[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5021_ as2650.r123\[0\]\[3\] as2650.r123_2\[0\]\[3\] _4008_ _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_79_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7216__A2 _2485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8413__A1 _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5227__A1 _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6293__I _1656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6972_ _1070_ _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6975__A1 _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5778__A2 _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8711_ _3344_ _3884_ _3313_ _3885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5923_ _1211_ _1302_ _1310_ _0058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_94_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8642_ as2650.stack\[4\]\[13\] _3819_ _3828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5854_ _1248_ _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4805_ _4212_ _4384_ _4385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8192__A3 _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8573_ _3764_ _3765_ _3766_ _3767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5785_ _1138_ _1181_ _1188_ _0042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_37_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8013__I _3247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7524_ _1615_ _2731_ _2772_ _2773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4736_ _4316_ _4317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7455_ _2702_ _2703_ _2704_ _2705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7152__A1 _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4667_ as2650.ins_reg\[4\] _4025_ as2650.ins_reg\[7\] _4248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_135_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6406_ _1744_ _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4505__A3 _4085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7386_ _1293_ _2639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4598_ _4178_ _4170_ _4179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6337_ _1642_ _1676_ _1692_ _1694_ _0088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9056_ _0217_ clknet_leaf_67_wb_clk_i as2650.r0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7455__A2 _2703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6268_ _0518_ _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7801__B _3042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8007_ _3223_ _3237_ _3241_ _3242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_9_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5219_ _0416_ _4414_ _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6199_ _1570_ _1571_ _1574_ _0070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8616__C _2620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7207__A2 _2455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8404__A1 _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7299__I _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6966__A1 _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5769__A2 _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8909_ _0070_ clknet_leaf_78_wb_clk_i as2650.ins_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8707__A2 _2550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4652__S _4010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7391__A1 _1843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4451__I as2650.cycle\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8882__CLK clknet_leaf_46_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8643__A1 _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7446__A2 _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6103__C1 _4393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8807__B _2530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6654__B1 _1972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4680__A2 _4092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4626__I _4206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_32_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6709__A1 _2003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5570_ _1001_ _1002_ _1003_ _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_102_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4521_ _4028_ _4102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8768__I _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7134__A1 _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7240_ _1777_ _2504_ _2506_ _2507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5145__B1 _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4452_ as2650.cycle\[0\] _4033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5696__A1 _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5696__B2 as2650.r123_2\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7171_ _2436_ _2442_ _2426_ _2443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_125_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6122_ _1506_ _1403_ _0604_ _1507_ _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_113_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_71_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6053_ _1439_ _1440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5004_ _4269_ _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_6_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7340__C _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8008__I _3242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6948__A1 as2650.r123_2\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6955_ as2650.r123_2\[0\]\[6\] _2223_ _2248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6412__A3 _1750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8452__B _3650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5620__A1 _4038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5906_ _1299_ _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6886_ _2185_ _2192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8625_ net40 _3713_ _3714_ _3817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5837_ _4214_ _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4806__S0 _4018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8556_ _3097_ _3750_ _3751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_22_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5923__A2 _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5768_ _1176_ _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7507_ _1354_ _2755_ _2756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4719_ _4068_ _4300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__7125__A1 _2393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8487_ _1696_ _3490_ _3684_ _2572_ _3685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__7582__I _2683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6700__B _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5699_ _1125_ _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7676__A2 _2692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7438_ _2687_ _2688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5687__A1 _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_49_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5687__B2 as2650.r123_2\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7369_ _2561_ _2625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9108_ _0269_ clknet_leaf_14_wb_clk_i net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8625__A1 net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7428__A2 _2677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5439__A1 _4017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9039_ _0200_ clknet_3_7_0_wb_clk_i as2650.pc\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6926__I _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6100__A2 _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4446__I _4026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6939__A1 _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7600__A2 _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5611__A1 _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5277__I _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5914__A2 _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_51_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7706__B _2950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9060__CLK clknet_leaf_39_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5142__A3 _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8616__A1 _3537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7419__A2 _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8616__B2 _3763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8092__A2 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7160__C _2431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6642__A3 _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4653__A2 _4233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5602__B2 _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6740_ _0537_ _1968_ _1838_ _2058_ _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6671_ _0751_ _0842_ _1992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7355__A1 _2591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5187__I _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7355__B2 _2611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8410_ _2899_ _0451_ _3610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5622_ _0351_ _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5905__A2 _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8341_ _3541_ _3542_ _3543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7107__A1 _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5553_ _0903_ _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_129_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4504_ _4079_ _4084_ _4085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8272_ _1398_ _2897_ _3476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5484_ _0921_ _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7223_ _1399_ _2490_ _2491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4435_ as2650.halted net10 _4016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7154_ _2392_ _2399_ _2425_ _2426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_119_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8447__B _3644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6105_ _1371_ _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7085_ _4317_ _1903_ _2364_ as2650.r123\[2\]\[0\] _2365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6094__A1 _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6036_ _4080_ _1229_ _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__7830__A2 _2861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4644__A2 _4072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5841__A1 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7987_ _2530_ _2406_ _3222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_42_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6938_ _0415_ _2219_ _2234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_74_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5097__I _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6869_ _2170_ _2180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8608_ _1122_ _3483_ _3800_ _3801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5357__C2 _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9083__CLK clknet_leaf_24_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8539_ _2252_ _3734_ _3735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__8201__I _3409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8074__A2 _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8920__CLK clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8076__C _2730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6085__A1 _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5832__A1 _4079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4635__A2 _4215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7487__I _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4904__I _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5060__A2 _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8837__A1 _2515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6312__A2 _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8065__A2 _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5470__I _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6076__A1 _4101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7812__A2 _2987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5823__A1 _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7910_ _3120_ _3124_ _3148_ _3149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8890_ _0051_ clknet_leaf_41_wb_clk_i as2650.psu\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7841_ as2650.pc\[9\] _3082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_110_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_52_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7772_ _3012_ _0898_ _3013_ _0912_ _3014_ _3015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4984_ _0426_ _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_23_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5051__A2 _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6723_ _2037_ _2042_ _2043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_71_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_20_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6654_ _0331_ _1966_ _1972_ _1974_ _1906_ _1975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_137_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5605_ _1027_ _1036_ _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6585_ _1906_ _1907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6551__A2 _4321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8324_ net53 net28 _3526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5536_ _0906_ _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8828__A1 _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8255_ _3458_ _3459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8943__CLK clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5467_ _0890_ _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7206_ _2457_ _2459_ _1563_ _2476_ _2477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_132_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8186_ _1648_ _3398_ _3405_ _3406_ _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5398_ _0759_ _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_28_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7137_ _2408_ _2272_ _2409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8056__A2 _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6067__A1 _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7803__A2 _3042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7068_ _1394_ _1449_ _2349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5814__A1 _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6019_ _0431_ _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_27_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7567__A1 _2592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5042__A2 _4304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7319__A1 _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6790__A2 _2069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_64_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_64_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_6_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4553__A1 _4017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8819__A1 _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6058__A1 _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7558__A1 _4391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5569__B1 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7010__I _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6230__A1 _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8770__A3 _3939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4570__S _4009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6533__A2 _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6370_ _1174_ _1048_ _1601_ _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_5321_ _0756_ _0757_ _0760_ _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6297__A1 _1592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8040_ _3268_ _4186_ _3270_ _3274_ _3275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_130_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5252_ _0691_ _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6836__A3 _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4847__A2 _4127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4809__I _4388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5183_ as2650.holding_reg\[5\] _0616_ _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6049__A1 _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8942_ _0103_ clknet_leaf_43_wb_clk_i as2650.stack\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_84_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7549__A1 _2796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8873_ _0034_ clknet_leaf_48_wb_clk_i as2650.stack\[6\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4544__I _4124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7824_ _3063_ _3065_ _3066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_97_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8761__A3 _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7755_ as2650.stack\[3\]\[6\] _1663_ _2999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4967_ _4331_ _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_75_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4783__A1 _4048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6706_ _2013_ _2025_ _2026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7686_ _1643_ _2930_ _2931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_4898_ as2650.r123\[1\]\[3\] as2650.r123\[0\]\[3\] as2650.r123_2\[1\]\[3\] as2650.r123_2\[0\]\[3\]
+ _4018_ _0339_ _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_137_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6637_ _1931_ _1958_ _1959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6524__A2 _4127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4535__A1 _4043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6568_ _0563_ _0765_ _1891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8307_ _4241_ _4271_ _3510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7804__B _3011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5519_ as2650.stack\[4\]\[9\] _0904_ _0918_ as2650.stack\[5\]\[9\] _0956_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6499_ _0353_ _1804_ _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6288__A1 _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8238_ _1207_ _3438_ _3444_ _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__9121__CLK clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4838__A2 _4188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8169_ as2650.stack\[6\]\[2\] _3393_ _3394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7788__A1 _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8354__C _3555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5263__A2 _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output30_I net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4454__I _4034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6212__A1 _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7260__I0 _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6212__B2 _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8989__CLK clknet_leaf_67_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6763__A2 _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7960__A1 _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7712__A1 as2650.stack\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7712__B2 as2650.stack\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8529__C _3687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7476__B1 _2690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4829__A2 _4374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4629__I _4209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_77_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8545__B _2629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6451__A1 _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5254__A2 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5870_ _0872_ _1244_ _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_61_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4821_ _4244_ _4400_ _4401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7951__A1 _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7540_ _1284_ _2536_ _2788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4752_ _4232_ _4234_ _4236_ _4332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__4765__A1 _4177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7471_ _2705_ _2720_ _2721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4683_ _4112_ _4263_ _4264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__5195__I as2650.holding_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7703__A1 _4095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4517__A1 _4089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6422_ _1629_ _1746_ _1757_ _0110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6353_ _1704_ _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5190__A1 _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5304_ _0659_ _0742_ _0743_ _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_66_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9072_ _0233_ clknet_leaf_41_wb_clk_i as2650.stack\[7\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6284_ _1648_ _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8023_ _1387_ _3258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5235_ _0652_ _0654_ _0675_ _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_130_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5493__A2 _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5166_ _0536_ _0606_ _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_111_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6037__A4 _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5097_ _0538_ _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8925_ _0086_ clknet_leaf_36_wb_clk_i as2650.stack\[4\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6993__A2 _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8856_ _0017_ clknet_leaf_55_wb_clk_i as2650.stack\[3\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8195__A1 as2650.stack\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_7807_ _3009_ _3048_ _3049_ _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7942__A1 as2650.addr_buff\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6745__A2 _2062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5999_ _0602_ _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8787_ _3937_ _3951_ _3956_ _3957_ _3958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4756__A1 as2650.holding_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7738_ _2446_ _2968_ _2981_ _1257_ _1317_ _2982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_71_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8498__A2 _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7669_ _2813_ _2906_ _2914_ _2470_ _2915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_123_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4771__A4 _4350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8422__A2 _3558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6028__A4 _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6433__A1 _1654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8084__C _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9017__CLK clknet_leaf_7_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4995__A1 _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8186__A1 _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7709__B _2946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7933__A1 _3089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4747__A1 _4326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6332__C _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5172__A1 _4370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5711__A3 _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7449__B1 _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_61_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_48_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5020_ _0284_ _0376_ _0377_ _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8275__B _2471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8413__A2 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5227__A2 _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6971_ _2261_ _1548_ _1567_ _2262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6975__A2 _4123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8710_ _1528_ _2522_ _3883_ _3884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_94_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5922_ as2650.stack\[0\]\[14\] _1300_ _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8177__A1 _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5853_ _1061_ _1246_ _1247_ _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_8641_ _1207_ _3821_ _3827_ _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_80_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7924__A1 _2813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4804_ as2650.r123\[2\]\[2\] as2650.r123_2\[2\]\[2\] _4011_ _4384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_22_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8572_ _3731_ _3733_ _2561_ _3766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_5784_ as2650.stack\[2\]\[13\] _1179_ _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4735_ _4315_ _4316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7523_ _2732_ _2734_ _2771_ _2727_ _2772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_120_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7454_ _0937_ _2265_ _2538_ _2704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_4666_ _4244_ _4247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6405_ _1174_ _1048_ _1591_ _1744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_7385_ _2531_ _2637_ _2638_ _2479_ _0192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4597_ _4066_ _4178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4910__A1 _4024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6336_ _1693_ _1680_ _1681_ _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8101__A1 _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_9055_ _0216_ clknet_leaf_65_wb_clk_i as2650.r0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6267_ _1629_ _1595_ _1634_ _0078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6112__B1 _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7455__A3 _2704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8006_ _2422_ _3240_ _3241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5218_ _0657_ _0569_ _0658_ _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7860__B1 _3087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6198_ _1572_ _1573_ _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8404__A2 _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5149_ _0589_ _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6415__A1 _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6966__A2 _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8908_ _0069_ clknet_leaf_78_wb_clk_i as2650.ins_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_60_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8707__A3 _2677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8839_ _0000_ clknet_leaf_1_wb_clk_i as2650.r123\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7915__A1 _2947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5828__I _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6718__A2 _2037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6194__A3 _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8140__S _3244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8340__A1 _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6103__B1 _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8643__A2 _3821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6103__C2 _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8807__C _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6654__A1 _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4968__A1 _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8542__C _3626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7906__A1 _3064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4642__I _4222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7953__I _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4520_ _4070_ _4100_ _4101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7134__A2 _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8331__A1 as2650.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4451_ as2650.cycle\[1\] _4032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5145__A1 _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7685__A3 _2833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6893__A1 _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7170_ _2438_ _2441_ _2442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6121_ as2650.psl\[5\] _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_112_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8634__A2 _3823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6052_ _4102_ _1438_ _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5003_ _0444_ _0445_ _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_26_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8398__A1 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6948__A2 _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7070__A1 _2344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6954_ _1034_ _2213_ _2221_ _2247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__8452__C _3294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5620__A2 _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5905_ _1044_ _1298_ _1084_ _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_74_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5648__I _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6885_ _1835_ _2186_ _2190_ _2191_ _0139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_74_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8024__I _2349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8624_ _1130_ _3558_ _3815_ _2485_ _3816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5836_ _0405_ _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8570__A1 _3063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5384__A1 _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8555_ _3062_ _3725_ _3727_ _3750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_5767_ _1175_ _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7506_ _2536_ _2749_ _2754_ _2755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_108_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4718_ _4298_ _4299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__7125__A2 _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8486_ _1360_ _3665_ _3683_ _3684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5698_ as2650.r123\[0\]\[3\] _1113_ _1124_ _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5136__A1 _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7437_ _2437_ _2687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4649_ _4229_ _4230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_107_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6884__A1 _4306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7368_ _2623_ _2563_ _2624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_9107_ _0268_ clknet_leaf_14_wb_clk_i net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8694__I _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6319_ _1671_ _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7428__A3 _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7299_ _0785_ _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5439__A2 _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7833__B1 _3072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9038_ _0199_ clknet_leaf_31_wb_clk_i as2650.pc\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4727__I _4307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8389__A1 _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6939__A2 _2213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7061__A1 _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5611__A2 _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8561__A1 _3602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5375__A1 _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7116__A2 _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5127__A1 _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6875__A1 _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5142__A4 _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7419__A3 _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6627__A1 _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6670_ _1895_ _1990_ _1950_ _1952_ _1991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_32_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5621_ _4288_ _1050_ _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5366__A1 _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8340_ _1404_ _0327_ _3542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5552_ as2650.stack\[3\]\[11\] _0948_ _0950_ _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7107__A2 _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4503_ _4080_ _4083_ _4084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8271_ _2606_ _2469_ _3475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5483_ _0909_ _0912_ _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7222_ _2489_ _2490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4434_ _4014_ _4015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_133_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7153_ _2402_ _2414_ _2420_ _2424_ _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__7632__B _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6618__A1 _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6104_ as2650.psu\[4\] _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_99_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7084_ _2363_ _2364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_98_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6094__A2 _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6035_ _1269_ _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5841__A2 _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7043__A1 _4195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7986_ _2268_ _4081_ _2393_ _3221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8791__A1 _3935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8872__CLK clknet_leaf_57_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6937_ _2228_ _2230_ _2233_ _0149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_74_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6868_ _2168_ _2179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8607_ _3797_ _3799_ _3800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7807__B _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5357__A1 _4222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5819_ _4307_ _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5357__B2 _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6799_ _2116_ _2117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8538_ _3731_ _3733_ _3734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6430__C _1744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5109__A1 _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8469_ _0725_ _0708_ _3667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_136_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6857__A1 _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6857__B2 as2650.stack\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7282__A1 _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4457__I _4037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6085__A2 _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5832__A2 _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5997__B _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7034__A1 _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8782__A1 _3951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8534__A1 _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5348__A1 _4221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4568__S _4009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6076__A2 _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8895__CLK clknet_leaf_51_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5823__A2 _4295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7025__A1 _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7840_ _3051_ _2686_ _3081_ _0204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_63_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8773__A1 _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5587__A1 _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7771_ as2650.stack\[0\]\[7\] _1192_ _2956_ as2650.stack\[1\]\[7\] _3014_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_51_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5198__I _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4983_ _0425_ _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_75_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6722_ _0592_ _0842_ _2042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8525__A1 _3326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5339__A1 _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6653_ _0334_ _1973_ _1918_ _1974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5604_ _0738_ _0871_ _0878_ _1035_ _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_20_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6584_ _4061_ _1811_ _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_8323_ _3479_ _3525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5535_ _0953_ _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8828__A2 _3952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8254_ _2391_ _3457_ _3458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5466_ _0903_ _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7205_ _2462_ _2475_ _2476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5397_ _0761_ _0768_ _0835_ _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_67_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8185_ _1696_ _3388_ _3385_ _3406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_101_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7136_ _2269_ _2408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6067__A2 _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7067_ _1253_ _1226_ _2314_ _2348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_100_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6018_ _1404_ _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5814__A2 _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6492__I _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9050__CLK clknet_leaf_64_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7969_ _1135_ _2731_ _2339_ _3206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7319__A2 _2576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7029__S _2294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5836__I _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5057__B _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4553__A2 _4133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_33_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_33_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_124_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6058__A2 _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7255__A1 _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_37_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5805__A2 _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8755__A1 _2257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7558__A2 _4233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6230__A2 _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8507__A1 _3021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4792__A2 _4371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5741__A1 _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5320_ _0758_ _0759_ _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_6_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7494__A1 _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5251_ _0396_ _0600_ _0690_ _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6297__A2 _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5182_ as2650.holding_reg\[5\] _0616_ _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6049__A2 _4296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8941_ _0102_ clknet_leaf_37_wb_clk_i as2650.stack\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9073__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8872_ _0033_ clknet_leaf_57_wb_clk_i as2650.stack\[6\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7201__I _2471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4480__A1 _4048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7549__A2 _2777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8746__A1 as2650.carry vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7823_ _3064_ _3034_ _2320_ _3065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_97_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8741__B _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7754_ as2650.stack\[7\]\[6\] _1297_ _2691_ as2650.stack\[6\]\[6\] _0914_ _2998_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_71_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4966_ _0391_ _0404_ _0408_ _0312_ _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6705_ _2023_ _2024_ _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4783__A2 _4055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7685_ _1688_ _1683_ _2833_ _2930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_4897_ _4213_ _0340_ _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4560__I _4140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8910__CLK clknet_leaf_9_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6636_ _1933_ _1957_ _1958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4535__A2 _4115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7871__I as2650.pc\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6567_ _1886_ _1889_ _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8306_ _3468_ _3509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5518_ as2650.stack\[2\]\[9\] _0952_ _0908_ as2650.stack\[1\]\[9\] _0954_ _0955_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_106_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6498_ _1820_ _1821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8237_ as2650.stack\[7\]\[12\] _3440_ _3444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_79_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5449_ _0886_ _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4838__A3 _4321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8168_ _3389_ _3393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7119_ _2258_ _2390_ _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8099_ _1490_ _3252_ _3329_ _0936_ _3330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_19_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_12_wb_clk_i_I clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4735__I _4315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8737__A1 _3904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output23_I net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7260__I1 _2522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6212__A2 _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7267__B _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4774__A2 _4353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5566__I _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4470__I as2650.cycle\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7712__A2 _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4526__A2 _4098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7714__C _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7476__A1 _1667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_51_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7476__B2 _2700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_26_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9096__CLK clknet_leaf_53_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8826__B _3990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7228__A1 _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6451__A2 _1750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8728__A1 _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8728__B2 _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8561__B _3755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7400__A1 _4128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7251__I1 _2515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4820_ _4238_ _4399_ _4400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7951__A2 _2842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5962__A1 _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4751_ _4178_ _4167_ _4331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5476__I _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4682_ _4261_ _4262_ _4263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7470_ _1598_ _2707_ _2719_ _1797_ _2720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7703__A2 _2416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6421_ _1632_ _1749_ _1752_ as2650.stack\[2\]\[3\] _1755_ _1757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__4517__A2 _4092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5714__A1 as2650.stack\[3\]\[13\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7624__C _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6352_ as2650.r123\[3\]\[3\] _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5303_ _0656_ _0674_ _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7467__A1 _4242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6283_ _0713_ _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_9071_ _0232_ clknet_leaf_42_wb_clk_i as2650.stack\[7\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8022_ _4322_ _3246_ _3256_ _3257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5234_ _0656_ _0659_ _0674_ _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XANTENNA__6690__A2 _2010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5165_ _4077_ _0426_ _0448_ _0583_ _4397_ _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_116_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5096_ net9 _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8027__I _4379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8924_ _0085_ clknet_leaf_30_wb_clk_i as2650.stack\[4\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8719__A1 _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6993__A3 _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8855_ _0016_ clknet_leaf_47_wb_clk_i as2650.stack\[3\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7806_ _2532_ _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8786_ _3951_ _3945_ _3937_ _3957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5998_ _1267_ _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7942__A2 _2803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7737_ _2979_ _2980_ _2981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4756__A2 _4332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4949_ _0387_ _4389_ _4337_ _4345_ _4334_ _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_71_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7668_ _2263_ _2913_ _2914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6619_ _4208_ _0369_ _1941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7599_ _2844_ _2845_ _2846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6130__A1 _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4692__A1 _4112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7630__A1 _2831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8956__CLK clknet_leaf_56_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6433__A2 _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8381__B _3534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8186__A2 _3398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5944__A1 as2650.psl\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4747__A2 _4113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7146__B1 _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7697__A1 _2940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5172__A2 _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7449__A1 as2650.stack\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7449__B2 as2650.stack\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7016__I _2293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4576__S _4154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4683__A1 _4112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6970_ _2260_ _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4435__A1 as2650.halted vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6975__A3 _2265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5921_ _1209_ _1302_ _1309_ _0057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_65_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8177__A2 _3398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8640_ as2650.stack\[4\]\[12\] _3823_ _3827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_94_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5852_ _4032_ _4118_ _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9111__CLK clknet_leaf_41_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7924__A2 _3146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4803_ _4382_ _4020_ _4383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8571_ _3725_ _3727_ _4092_ _3765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5935__A1 _4156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5783_ _1133_ _1181_ _1187_ _0041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7522_ _2759_ _2769_ _2770_ _2771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4734_ _4309_ _4314_ _4315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7453_ _1596_ _4062_ _2703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4665_ _4245_ _4246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6404_ _1654_ _1712_ _1743_ _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_128_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7384_ _2633_ _2634_ _4050_ _2638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4596_ as2650.psl\[3\] as2650.carry _4177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6335_ _1645_ _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_1_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4910__A2 _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8101__A2 _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9054_ _0215_ clknet_leaf_64_wb_clk_i as2650.r0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6112__A1 _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6266_ _1632_ _1604_ _1594_ _1633_ _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__6112__B2 _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8005_ _1345_ _1455_ _3239_ _2656_ _3240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__7860__A1 _2947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5217_ _0469_ _0568_ _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8979__CLK clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7860__B2 _2599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6197_ _1564_ _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5148_ _0588_ _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7612__A1 _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5079_ _4019_ _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_71_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8907_ _0068_ clknet_leaf_74_wb_clk_i as2650.r123_2\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7596__I _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6179__A1 _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8838_ _3999_ _4000_ _3049_ _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_38_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7915__A2 _3150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5926__A1 _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8769_ _3940_ _3938_ _3941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7679__A1 _2689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7679__B2 _2915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8340__A2 _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6103__A1 _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6654__A2 _1966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7603__A1 _2843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8823__C _3659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4968__A2 _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5090__A1 _4213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6590__A1 _4400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8331__A2 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4450_ _4028_ _4030_ _4031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6893__A2 _2012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6120_ as2650.overflow _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_124_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6051_ _1246_ _1247_ _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4656__A1 _4232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5002_ _0319_ _0301_ _0399_ _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_61_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6953_ _1028_ _2219_ _2246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4959__A2 _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5904_ _1297_ _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_81_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6884_ _4306_ _4322_ _2071_ _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_39_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8623_ _3519_ _3808_ _3811_ _3814_ _2481_ _3815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_62_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5835_ _1229_ _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8570__A2 _2296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8554_ _2296_ _3748_ _3749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_124_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5384__A2 _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5766_ _0895_ as2650.psu\[1\] _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7505_ _2445_ _2733_ _2753_ _2754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4717_ _4297_ _4298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8485_ _3666_ _3680_ _3682_ _3500_ _3473_ _3683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__5664__I _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5697_ _1123_ _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_135_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7436_ _2685_ _2686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5136__A2 _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4648_ as2650.r0\[1\] _4229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6333__A1 _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__9007__CLK clknet_leaf_76_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6884__A2 _4322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7367_ _2622_ _2623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_122_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4579_ _4152_ _4160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_9106_ _0267_ clknet_leaf_13_wb_clk_i net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8086__A1 _3303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6318_ _1623_ _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_46_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7298_ _2480_ _2556_ _2557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_81_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7833__A1 _2793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6636__A2 _1957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9037_ _0198_ clknet_leaf_30_wb_clk_i as2650.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6249_ _1611_ _1595_ _1618_ _0076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_89_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_18_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7061__A2 _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_58_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_58_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_73_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5072__A1 _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8561__A2 _3747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6572__A1 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5375__A2 _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5127__A2 _4319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4886__A1 _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4886__B2 _4371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8077__A1 _3271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7419__A4 _2668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7824__A1 _3063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7588__B1 _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5063__A1 _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7169__C _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8001__A1 _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5620_ _4038_ _1049_ _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5551_ as2650.r123\[0\]\[3\] _0878_ _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4602__B _4165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8304__A2 _3506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4502_ _4082_ _4083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8270_ _3447_ _3463_ _3471_ _3472_ _3473_ _3474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5482_ _0898_ _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7913__B _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7221_ _0937_ _2489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4433_ _4013_ _4014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4877__A1 _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7152_ _1050_ _2423_ _2424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6079__B1 _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6103_ _1487_ _1488_ _0605_ _1213_ _4393_ _0897_ _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_115_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7083_ _0940_ _4315_ _2362_ _2363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_59_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6034_ _4049_ _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8744__B _3916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7043__A2 _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8240__A1 _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7985_ _2640_ _3220_ _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5659__I _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8035__I _3269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6936_ _0981_ _2231_ _2221_ _2232_ _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_78_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6867_ _2166_ _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8606_ _1122_ _3525_ _3798_ _2668_ _2437_ _3799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_50_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5818_ as2650.psu\[5\] _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5357__A2 _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6798_ _2114_ _2115_ _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_8537_ _4365_ _3732_ _3733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5749_ as2650.stack\[6\]\[8\] _1164_ _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5109__A2 _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8468_ _3463_ _3661_ _3517_ _3666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_68_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7823__B _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7419_ _1845_ _2281_ _2288_ _2668_ _2669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
X_8399_ _2845_ _3582_ _3599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8059__A1 _3258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7542__C _2789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8059__B2 _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5343__B _4174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4738__I _4318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7282__A2 _4122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5293__A1 _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7034__A2 _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5045__A1 as2650.holding_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8782__A2 _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8534__A2 _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8298__A1 _2712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6848__A2 _2069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7733__B _2894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4648__I as2650.r0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5823__A3 _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7025__A2 _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8773__A2 _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7770_ as2650.stack\[3\]\[7\] _1663_ _3013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6784__A1 _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4982_ _0424_ _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6721_ _4208_ _1951_ _2041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_leaf_3_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_60_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6652_ _0883_ _4116_ _1811_ _1973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__5339__A2 _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5603_ _1028_ _0882_ _0889_ _1034_ _0930_ _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_6583_ _1800_ _1905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8322_ _3489_ _3522_ _3524_ _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8289__A1 _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5534_ as2650.stack\[2\]\[10\] _0969_ _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8739__B _3303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8253_ _2399_ _3453_ _3456_ _3457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_118_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5465_ _0895_ _0902_ _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8458__C _3656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7204_ _2336_ _1348_ _2463_ _2468_ _2474_ _2475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
X_8184_ as2650.stack\[6\]\[6\] _3390_ _3405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5396_ _0562_ _0762_ _0767_ _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_82_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7135_ _2268_ _1334_ _2257_ _2343_ _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_113_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4558__I _4135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6067__A3 _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7066_ _2316_ _2344_ _2322_ _2346_ _2347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_28_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8474__B _3671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6017_ _1403_ _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8213__A1 _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8764__A2 _3935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7968_ _2591_ _3203_ _3204_ _2685_ _3205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6919_ _1834_ _2208_ _2217_ _0147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_74_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7899_ _3110_ _3138_ _3049_ _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_70_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7319__A3 _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6527__A1 _1837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6013__I _4392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5750__A2 _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_41_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4468__I _4043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_73_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_73_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__8452__A1 _3626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7255__A2 _2517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5266__A1 _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8204__A1 _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6215__B1 _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5569__A2 _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5033__A4 _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7715__B1 _2958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_80_wb_clk_i_I clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7019__I as2650.addr_buff\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5741__A2 _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8691__A1 _3851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7494__A2 _2416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5250_ _0689_ _0396_ _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8862__CLK clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4701__B1 _4279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5181_ _0486_ _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8443__A1 _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6049__A3 _4331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5257__A1 _4172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8940_ _0101_ clknet_leaf_42_wb_clk_i as2650.stack\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8871_ _0032_ clknet_leaf_54_wb_clk_i as2650.stack\[6\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_37_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4480__A2 _4049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8746__A2 _3916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7822_ _0784_ _4215_ _3064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7753_ as2650.stack\[4\]\[6\] _2836_ _1176_ as2650.stack\[5\]\[6\] _2997_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4965_ _0405_ _0407_ _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6704_ _0413_ _1965_ _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7684_ _1693_ _2878_ _2929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4896_ as2650.r123\[2\]\[3\] as2650.r123_2\[2\]\[3\] _0339_ _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5980__A2 _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6635_ _1938_ _1956_ _1957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7182__A1 _4054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6524__A4 _1846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6566_ _1887_ _1888_ _1889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5732__A2 _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4535__A3 _4075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8305_ _3465_ _3503_ _3504_ _3507_ _3508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_69_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5517_ as2650.stack\[0\]\[9\] _0953_ _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_118_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6497_ _4225_ _1812_ _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8236_ _1205_ _3437_ _3443_ _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8682__A1 _3838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5448_ _0885_ _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4838__A4 _4417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8167_ _1721_ _3386_ _3392_ _0220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_114_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5379_ _0817_ _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_99_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8434__A1 _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7118_ _2136_ _0787_ _2386_ _2389_ _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_8098_ _4286_ _3251_ _3329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5248__A1 _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7049_ _1474_ _1249_ _2331_ _2332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_74_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6996__A1 _4091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6008__I _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_8_wb_clk_i_I clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output16_I net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5847__I _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_15_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7173__A1 _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8885__CLK clknet_leaf_52_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6920__A1 _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4526__A3 _4106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8379__B _3579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8122__B1 _3350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7476__A2 _2689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8425__A1 _3595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7228__A2 _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4926__I _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6987__A1 _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6451__A3 _1766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8728__A2 _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6739__A1 _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8561__C _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7400__A2 _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4661__I _4241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7177__C _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4750_ _4325_ _4329_ _4330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5962__A2 _4376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4681_ _4093_ _4096_ _4262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6420_ _1620_ _1746_ _1756_ _0109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4517__A3 _4097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5714__A2 _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6351_ _1703_ _0093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5302_ _0656_ _0674_ _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9070_ _0231_ clknet_leaf_41_wb_clk_i as2650.stack\[7\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7467__A2 _2716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6282_ _1642_ _1637_ _1647_ _0080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8021_ _3250_ _3254_ _3246_ _3255_ _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7921__B _2735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5233_ _0663_ _0673_ _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_88_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7219__A2 _2484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5164_ _0604_ _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_69_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4836__I _4415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7212__I _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5095_ _0536_ _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8923_ _0084_ clknet_leaf_32_wb_clk_i as2650.stack\[4\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5650__A1 _4142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8719__A2 _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6993__A4 _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8854_ _0015_ clknet_leaf_68_wb_clk_i as2650.r123\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_52_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7805_ _2831_ _3045_ _3047_ _2829_ _3048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XPHY_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8785_ _2505_ _3952_ _3955_ _1279_ _3956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_5997_ _1367_ _1382_ _1383_ _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8043__I _2622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7736_ _1374_ _2851_ _2980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4948_ _0385_ _0390_ _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7667_ _2909_ _2912_ _2913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4879_ _4232_ _4234_ _4236_ _4153_ _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_4
XFILLER_138_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6618_ _1890_ _1897_ _1939_ _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7598_ _1630_ net8 _2845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6902__A1 _2147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6549_ _0828_ _0854_ _1872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8104__B1 _3333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8219_ as2650.stack\[7\]\[6\] _3424_ _3431_ _3408_ _3432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_121_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8407__A1 _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4692__A2 _4061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4746__I as2650.holding_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5641__A1 _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6961__I as2650.addr_buff\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7146__A1 _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7146__B2 _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7697__A2 _2904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5526__B _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9063__CLK clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_3_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6201__I _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7449__A2 _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4683__A2 _4263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8572__B _2561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5632__A1 _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4435__A2 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5920_ as2650.stack\[0\]\[13\] _1300_ _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5851_ _1058_ _1053_ _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__7385__A1 _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4802_ _4381_ _4382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_94_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8570_ _3063_ _2296_ _3764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5782_ as2650.stack\[2\]\[12\] _1183_ _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_128_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7521_ _2460_ _2770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4733_ _4313_ _4314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7452_ _1597_ _1577_ _2702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7688__A2 net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4664_ _4244_ _4245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6403_ _1741_ _1717_ _1710_ _1742_ _1743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_7383_ _2613_ _2636_ _2637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4595_ _4175_ _4158_ _4176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_9122_ _0283_ clknet_leaf_44_wb_clk_i as2650.psu\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6334_ as2650.stack\[4\]\[5\] _1677_ _1692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9053_ _0214_ clknet_leaf_70_wb_clk_i as2650.r0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6265_ as2650.stack\[5\]\[3\] _1616_ _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_142_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6112__A2 _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8004_ _4079_ _1433_ _3238_ _3239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5216_ _0469_ _0568_ _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7860__A2 _3092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6196_ _1401_ _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4674__A2 _4224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8038__I _2898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4566__I _4146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5147_ _0533_ _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7612__A2 _2858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5078_ as2650.r123_2\[1\]\[5\] _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_72_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8482__B _3579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8906_ _0067_ clknet_leaf_62_wb_clk_i as2650.r123_2\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_53_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8837_ _2515_ _3997_ _4000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7376__A1 _2591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6179__A2 _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8768_ _1261_ _3940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__9086__CLK clknet_leaf_25_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7128__A1 _4301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7719_ _2780_ _2937_ _2791_ _2964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8699_ _1432_ _3872_ _3873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_138_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5065__C _4165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5860__I _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8923__CLK clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6103__A2 _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7603__A2 _2849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5090__A2 _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5917__A2 _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7119__A1 _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6590__A2 _1911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7027__I _4093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8619__A1 _3626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6866__I _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6050_ _4038_ _1436_ _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_input7_I io_in[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5001_ _0319_ _0324_ _0398_ _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_113_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_22_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6952_ _2242_ _2243_ _2245_ _0152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7070__A3 _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5903_ _1296_ _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7358__A1 _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6883_ as2650.r123_2\[1\]\[0\] _2189_ _2190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6106__I net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8622_ _1130_ _3480_ _3813_ _3654_ _3175_ _3814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_5834_ _1073_ _4087_ _4144_ _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_126_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8553_ _3062_ _3731_ _3733_ _3748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_10_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5765_ _1173_ _1174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6581__A2 _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7504_ _2710_ _2749_ _2752_ _2263_ _2753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4716_ _4166_ _4069_ _4297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8484_ _2970_ _3681_ _3682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_120_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5696_ _1122_ _1089_ _1097_ as2650.r123_2\[0\]\[3\] _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_124_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7435_ _2684_ _2685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4647_ _4227_ _4228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7530__A1 _2539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8946__CLK clknet_leaf_33_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6333__A2 _1662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7366_ _2255_ _2622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6884__A3 _2071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4578_ _4158_ _4159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9105_ _0266_ clknet_leaf_13_wb_clk_i net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6317_ as2650.stack\[4\]\[2\] _1677_ _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8908__D _0069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8086__A2 _2014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7297_ _2537_ _2544_ _2555_ _2431_ _2556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6097__A1 _4006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9036_ _0197_ clknet_leaf_40_wb_clk_i as2650.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7833__A2 _3070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6248_ _1615_ _1604_ _1594_ _1617_ _1618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_83_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5844__A1 _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6179_ _1544_ _1549_ _1555_ _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7597__A1 _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_opt_3_0_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5072__A2 _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6016__I _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6021__A1 _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6572__A2 _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4886__A2 _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8077__A2 _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7285__B1 _2541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__9101__CLK clknet_leaf_13_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7588__A1 as2650.stack\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7588__B2 as2650.stack\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5599__B1 _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5063__A2 _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6563__A2 _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5765__I _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5550_ _0964_ _0985_ _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4574__A1 as2650.holding_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4501_ _4034_ _4081_ _4082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5481_ as2650.stack\[4\]\[8\] _0904_ _0918_ as2650.stack\[5\]\[8\] _0919_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_144_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7512__A1 as2650.stack\[4\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7220_ _4189_ _1317_ _2488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4432_ _4012_ _4013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_126_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4877__A2 _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7151_ _2343_ _2422_ _2423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6079__A1 _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6102_ _0783_ _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_28_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6079__B2 _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7082_ _2359_ _2362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6033_ _4292_ _1227_ _1419_ _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7579__A1 _2777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7579__B2 _2732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8316__I _3473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7043__A3 _2325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8240__A2 _3438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7984_ as2650.pc\[14\] _2731_ _3219_ _3220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6935_ _0980_ _2219_ _2232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8760__B _2883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_63_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6866_ _1635_ _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6003__A1 _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7376__B _2631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8605_ _2862_ _3792_ _3151_ _3798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5817_ _1211_ _1198_ _1212_ _0050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6797_ _4210_ _2036_ _2042_ _2115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_10_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4565__A1 _4142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8536_ _1488_ _0796_ _3732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5748_ _1162_ _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8467_ _1650_ _3491_ _3664_ _3498_ _3665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7503__A1 _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5679_ _1107_ _1099_ _1100_ _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA_clkbuf_leaf_31_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7418_ _1417_ _4081_ _1545_ _2668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_8398_ net32 _3597_ _3598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_117_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7349_ _1439_ _2606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8059__A2 _2651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5817__A1 _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9019_ _0180_ clknet_leaf_8_wb_clk_i as2650.holding_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5293__A2 _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8226__I _3436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8231__A2 _3440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7990__A1 _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_70_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7742__A1 _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4556__A1 _4007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4859__A2 _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4929__I _4375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6481__A1 _4131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4664__I _4244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4981_ _0419_ _0421_ _0423_ _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_2
X_6720_ _2038_ _2039_ _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6651_ _1387_ _1839_ _1970_ _1971_ _1972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5495__I as2650.r123\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7733__A1 _2882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5602_ _1029_ _1030_ _1033_ _0957_ _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_34_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6582_ _1835_ _1852_ _1866_ _1904_ _0123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_118_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8321_ net29 _3523_ _3191_ _3524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5533_ _0899_ _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8289__A2 _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8252_ _3454_ _3455_ _1334_ _2883_ _3456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_121_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5464_ as2650.psu\[1\] _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7203_ _1523_ _2470_ _2473_ _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8183_ _1734_ _3398_ _3403_ _3404_ _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5395_ _0832_ _0833_ _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7215__I _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7134_ _1426_ _2405_ _2406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7065_ _1272_ _2345_ _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8474__C _2622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6016_ _1402_ _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_74_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7967_ _2462_ _2782_ _3194_ _3204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7972__A1 as2650.pc\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4786__A1 _4362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6918_ _2210_ _2211_ _2216_ _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7818__C _2789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7898_ _2831_ _3135_ _3137_ _2829_ _3138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7319__A4 _2574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7724__A1 _1738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6849_ _2013_ _2151_ _2163_ _1852_ _2164_ _0130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_11_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8519_ _3489_ _3712_ _3715_ _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_108_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5354__B _4258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4749__I _4328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6964__I _4092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8452__A2 _3629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5266__A2 _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_46_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4484__I _4064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8204__A2 _3419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6215__A1 _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5018__A2 _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6215__B2 _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_42_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_42_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_3275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7963__A1 _2537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6518__A2 _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4659__I _4203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8691__A2 _3866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6079__C _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4701__A1 _4259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5180_ _4135_ _0620_ _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8870_ _0031_ clknet_leaf_57_wb_clk_i as2650.stack\[6\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_97_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7403__B1 _2653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4480__A3 _4056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7821_ _3062_ _3063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7954__A1 _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4768__A1 _4140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4964_ _0395_ _4191_ _0406_ _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_7752_ _2760_ _2996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_75_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6703_ _2021_ _2022_ _2023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_71_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7706__A1 _2947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7683_ _2830_ _2926_ _2928_ _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4895_ _4011_ _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_71_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6114__I _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6634_ _1940_ _1955_ _1956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7182__A2 _4122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5193__A1 _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6565_ _4229_ _0839_ _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5953__I _4223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8304_ _2625_ _3506_ _3507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5516_ _0903_ _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6496_ _1818_ _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8131__A1 _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8235_ as2650.stack\[7\]\[11\] _3440_ _3443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5447_ _4311_ _0884_ _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8682__A2 _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7890__B1 _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5378_ _0795_ _0798_ _0816_ _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_8166_ _1614_ _3388_ _3390_ as2650.stack\[6\]\[1\] _3384_ _3392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_120_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7117_ _0436_ _0543_ _0607_ _2388_ _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_141_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8097_ _3323_ _3325_ _3270_ _3327_ _3328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_86_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7048_ _2330_ _2331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6996__A2 _2286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7945__A1 _2947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8999_ _0160_ clknet_leaf_10_wb_clk_i as2650.addr_buff\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4759__A1 _4162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6452__C _1773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5420__A2 _4304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6024__I _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7173__A2 _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5184__A1 _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5863__I _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6920__A2 _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8122__A1 _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8122__B2 _3351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4479__I _4059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8673__A2 _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6694__I _4390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7228__A3 _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6436__A1 _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6987__A2 _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4942__I _4335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5259__B _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5962__A3 _4188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4680_ _4260_ _4092_ _4261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_109_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_30_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7164__A2 _2432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6869__I _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6350_ as2650.r123\[3\]\[2\] _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4922__A1 _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5301_ _0654_ _0739_ _0740_ _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6281_ _1646_ _1625_ _1607_ as2650.stack\[5\]\[5\] _1593_ _1647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__6124__B1 _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8664__A2 _3846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5232_ _0664_ _0668_ _0672_ _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_8020_ _0880_ _2700_ _3255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5163_ _0603_ _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6427__A1 _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7624__B1 _2867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5094_ _0535_ _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8922_ _0083_ clknet_leaf_36_wb_clk_i as2650.stack\[4\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6109__I _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5650__A2 _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7649__B _2894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8853_ _0014_ clknet_leaf_65_wb_clk_i as2650.r123\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7927__A1 _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5948__I _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7804_ _2438_ _3046_ _3011_ _3047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_8784_ _2428_ _0881_ _3954_ _3955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XPHY_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5996_ _4072_ _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7735_ _4094_ _2809_ _2979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_33_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4947_ _0386_ _0389_ _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_123_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7666_ _2910_ _2911_ _1335_ _2912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4878_ _4356_ _0318_ _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6617_ _1893_ _1896_ _1939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5166__A1 _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7597_ _1630_ _0429_ _2844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__6902__A2 _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4913__A1 _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6548_ _1870_ _0822_ _1871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8104__A1 _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6115__B1 _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6479_ _0291_ _1095_ _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8218_ _1738_ _3412_ _3431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_82_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8407__A2 _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8149_ _1527_ _3376_ _3377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6019__I _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5641__A2 _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8852__CLK clknet_leaf_68_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7933__A4 _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4601__B1 _4172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8343__A1 _3540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7146__A2 _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5157__A1 _4218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7313__I _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6409__A1 _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5632__A2 _4121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7469__B _2718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_93_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7909__A1 as2650.pc\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5768__I _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4840__B1 _4417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5850_ _1244_ _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7385__A2 _2637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4801_ as2650.r0\[2\] _4381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5396__A1 _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5781_ _1126_ _1180_ _1186_ _0040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_72_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7520_ _2760_ _2734_ _2768_ _2769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_72_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4732_ _4311_ _4312_ _4313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7137__A2 _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7451_ _2469_ _2701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4663_ _4023_ _4106_ _4244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6896__A1 _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6402_ as2650.stack\[3\]\[7\] _1714_ _1742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_7382_ _4050_ _2633_ _2636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4594_ _4174_ _4175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_9121_ _0282_ clknet_leaf_45_wb_clk_i as2650.psu\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6333_ _1636_ _1662_ _1691_ _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8637__A2 _3820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6648__A1 _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9052_ _0213_ clknet_leaf_66_wb_clk_i as2650.r0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6264_ _1631_ _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8003_ _1271_ _1352_ _0352_ _3238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5215_ _0655_ _0570_ _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6195_ _0945_ _1557_ _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5146_ _0586_ _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8270__B1 _3471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5077_ _4012_ as2650.r123\[1\]\[5\] _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_42_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8875__CLK clknet_leaf_46_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6820__A1 _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8905_ _0066_ clknet_leaf_62_wb_clk_i as2650.r123_2\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5678__I as2650.r123\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4582__I _4140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8836_ _2514_ _3992_ as2650.psu\[3\] _3999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7376__A2 _2619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5387__A1 _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8767_ _0334_ _1092_ _3939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5979_ _1365_ _0602_ _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_55_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7718_ _2937_ _2954_ _2960_ _2961_ _2962_ _2963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_40_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8325__A1 net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7128__A2 _4084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8698_ _2658_ _1461_ _2400_ _3871_ _3872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__5139__A1 _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7649_ _2882_ _2893_ _2894_ _2895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_126_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6302__I _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7064__A1 _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6972__I _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4492__I _4063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8564__A1 _3093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9030__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7119__A2 _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6878__A1 _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__8619__A2 _3810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5000_ _4270_ _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8898__CLK clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4656__A3 _4236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_85_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7055__A1 _2334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_opt_3_1_wb_clk_i clknet_opt_3_0_wb_clk_i clknet_opt_3_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_93_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6951_ _1022_ _2231_ _2214_ _2244_ _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_81_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5498__I _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5902_ _0911_ _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6882_ _2188_ _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7358__A2 _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8555__A1 _3062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_8621_ _3180_ _3812_ _3813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5369__A1 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5833_ _1214_ _1221_ _1227_ _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_34_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8552_ _3088_ _3746_ _3747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_124_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8307__A1 _4241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5764_ _1043_ _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7503_ _1439_ _2750_ _2751_ _2752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4715_ _4131_ _4295_ _4296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
X_8483_ _2932_ _3627_ _2973_ _3681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7515__C1 as2650.stack\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5695_ _1121_ _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7434_ _2683_ _2684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_129_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4646_ _4226_ _4227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7530__A2 _2706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7365_ _2439_ _2620_ _2621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4577_ _4156_ _4157_ _4158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5961__I _4294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9104_ _0265_ clknet_leaf_13_wb_clk_i net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6316_ _1672_ _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7296_ _2553_ _2554_ _2555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_103_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7294__A1 _2547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6097__A2 _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8049__I _3247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9035_ _0196_ clknet_leaf_40_wb_clk_i as2650.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7294__B2 _2552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6247_ as2650.stack\[5\]\[1\] _1616_ _1617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_103_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6178_ _1550_ _1551_ _1552_ _1554_ _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__8493__B _3572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7046__A1 _2314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5129_ _0562_ _0567_ _0570_ _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_131_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7597__A2 _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8794__A1 _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_129_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8819_ _2533_ _3985_ _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_81_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6021__A2 _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5780__A1 as2650.stack\[2\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_67_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_67_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_138_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5871__I _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7285__A1 _2434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8785__A1 _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8537__A1 _4365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4574__A2 _4154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4500_ _4053_ _4031_ _4081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5480_ _0907_ _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4431_ _4011_ _4012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5523__A1 _4377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5523__B2 _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7150_ _4049_ _1270_ _2421_ _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_99_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6079__A2 _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6101_ as2650.psu\[7\] _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_98_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7276__A1 _2334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7081_ _2360_ _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5826__A2 _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6032_ _4145_ _0927_ _1418_ _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9076__CLK clknet_leaf_53_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8776__A1 _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7983_ _3209_ _3218_ _2727_ _3219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_78_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6934_ _2218_ _2231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8528__A1 _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6865_ _1727_ _2167_ _2176_ _0134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_126_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5956__I _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7200__A1 _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6003__A2 _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8913__CLK clknet_leaf_9_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8604_ _2892_ _3150_ _3797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4860__I _4332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5816_ as2650.stack\[1\]\[14\] _1196_ _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6796_ _0710_ _2076_ _2114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8535_ _3673_ _3676_ _3730_ _3693_ _3731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_5747_ _1162_ _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4565__A2 _4145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8466_ _3663_ _3664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8488__B _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5678_ as2650.r123\[0\]\[1\] _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_136_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7503__A2 _2750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8700__A1 _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7417_ _1240_ _1433_ _2380_ _2667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4629_ _4209_ _4210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8397_ _3562_ _3563_ _3597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7348_ _1430_ _2319_ _2605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7267__A1 _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7279_ _2382_ _2390_ _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_49_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5817__A2 _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9018_ _0179_ clknet_leaf_7_wb_clk_i as2650.holding_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8767__A1 _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output39_I net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7990__A2 _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5866__I _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7742__A2 _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4556__A2 _4136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5753__A1 _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7258__A1 _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5808__A2 _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7321__I _2574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8758__A1 _2530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7430__A1 _2311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4980_ _4218_ _0422_ _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_64_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7981__A2 _3215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5992__A1 _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6650_ _1815_ _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5601_ as2650.stack\[3\]\[14\] _0893_ _0900_ as2650.stack\[2\]\[14\] _1032_ _1033_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_73_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5744__A1 _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6581_ _1867_ _1903_ _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8320_ _3459_ _3523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5532_ as2650.stack\[3\]\[10\] _0967_ _0950_ _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7497__A1 _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8251_ _2311_ _1442_ _2416_ _3455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5463_ as2650.stack\[3\]\[8\] _0893_ _0900_ as2650.stack\[2\]\[8\] _0901_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_117_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7202_ _2472_ _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8182_ _1693_ _3395_ _3396_ _3404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_132_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5394_ as2650.r0\[7\] _4318_ _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7249__A1 _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7133_ _2286_ _2404_ _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7064_ _1450_ _2343_ _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6015_ net7 _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6472__A2 _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4855__I _4165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8749__A1 _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8771__B _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7421__A1 _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7966_ _1021_ _2961_ _3194_ _2996_ _3202_ _3203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7972__A2 _3207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6917_ _1589_ _2213_ _2215_ _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4786__A2 _4364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5686__I as2650.pc\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7897_ _3113_ _3136_ _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_126_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4590__I _4170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6848_ as2650.r123_2\[2\]\[7\] _2069_ _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_10_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5735__A1 _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6779_ _0607_ _1853_ _2097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8518_ net35 _3713_ _3714_ _3715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7488__A1 _2735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8449_ _1282_ _3571_ _3645_ _3647_ _2255_ _3648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_87_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6310__I _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8959__CLK clknet_leaf_47_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7660__A1 _2898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6215__A2 _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7412__A1 _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7412__B2 _2662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4777__A2 _4356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5974__A1 _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5596__I _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7715__A2 _2957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_11_wb_clk_i clknet_3_2_0_wb_clk_i clknet_leaf_11_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_122_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7479__A1 _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7100__B1 _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7403__A1 _2647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7820_ as2650.addr_buff\[0\] _3062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4480__A4 _4060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6823__C _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7751_ _2983_ _2994_ _2995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4768__A2 _4168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4963_ _4190_ _0399_ _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6702_ _0458_ _1808_ _1802_ _2022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7682_ _1640_ _2878_ _2927_ _2928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5439__C _4285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4894_ _0337_ _4020_ _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7706__A2 _2935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6633_ _1945_ _1954_ _1955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6564_ _0751_ _0465_ _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8303_ _4090_ _3505_ _3506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5515_ _0898_ _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_121_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6495_ _1817_ _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7226__I _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4940__A2 _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8234_ _1203_ _3437_ _3442_ _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_69_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5446_ _4140_ _0874_ _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_86_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7890__A1 _2843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8165_ _1709_ _3386_ _3391_ _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7890__B2 _2796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5377_ _4139_ _0804_ _0815_ _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__8485__C _3473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7116_ _2387_ _0357_ _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8096_ _3326_ _0510_ _3327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7047_ _4089_ _2283_ _2330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4456__A1 _4031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8998_ _0159_ clknet_3_3_0_wb_clk_i as2650.addr_buff\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_70_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7945__A2 _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7949_ _2813_ _3179_ _3183_ _3186_ _3187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8520__I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5184__A2 _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6381__A1 _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6040__I _4031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8122__A2 _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7580__B _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7633__A1 _2830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6436__A2 _1766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6924__B _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8189__A2 _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7936__A2 _3173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4922__A2 _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5300_ _0652_ _0675_ _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6124__A1 _4173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6280_ _1645_ _1646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6124__B2 _4207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5231_ _0670_ _0671_ _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_9_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5162_ net1 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7624__A1 _2857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6427__A2 _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7624__B2 _2870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5093_ _0530_ _0532_ _0534_ _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_111_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8921_ _0082_ clknet_leaf_33_wb_clk_i as2650.stack\[5\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5650__A3 _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8852_ _0013_ clknet_leaf_68_wb_clk_i as2650.r123\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7927__A2 _2686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7803_ _2779_ _3042_ _3043_ _3046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_64_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5938__A1 _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8783_ _1610_ _3940_ _3953_ _3954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5995_ _1285_ _1378_ _1380_ _1381_ _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6125__I as2650.psl\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7734_ _2843_ _2975_ _2978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5169__C _4204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4946_ _0297_ _0306_ _0303_ _0388_ _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_127_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7665_ as2650.addr_buff\[4\] _2285_ _2598_ _2881_ _2890_ _2710_ _2911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai222_1
X_4877_ _0318_ _0320_ _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6616_ _1934_ _1937_ _1889_ _1886_ _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__6363__A1 _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7596_ _1052_ _2843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6547_ _0747_ _0829_ _1870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8104__A2 _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6115__A1 _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6478_ _1800_ _1801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6115__B2 _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8217_ _1734_ _3410_ _3429_ _3430_ _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_134_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5429_ _0862_ _0863_ _0866_ _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_0_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8148_ _2076_ _2377_ _3375_ _3376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8079_ _3268_ _3309_ _3310_ _3311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_48_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7918__A2 _3141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output21_I net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5929__A1 _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6035__I _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4601__A1 _4171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7146__A3 _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5157__A2 _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7854__A1 _3063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7606__A1 _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6409__A2 _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5093__A1 _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4953__I _4115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5632__A3 _4119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4840__A1 _4377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7909__A2 _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4840__B2 _4189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8031__A1 _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4800_ _4203_ _4380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5396__A2 _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5780_ as2650.stack\[2\]\[11\] _1183_ _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6593__A1 _4379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4731_ _4297_ _4300_ _4312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8334__A2 _3535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7450_ _2693_ _2696_ _2698_ _2699_ _2700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__6345__A1 _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4662_ _4242_ _4243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_11_wb_clk_i_I clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7542__B1 _2787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6401_ _1656_ _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6896__A2 _2012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7381_ _2633_ _2634_ _2635_ _0191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_134_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4593_ as2650.psl\[3\] _4173_ _4174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9120_ _0281_ clknet_3_6_0_wb_clk_i net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8098__A1 _4286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6332_ as2650.stack\[4\]\[4\] _1665_ _1690_ _1660_ _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_9051_ _0212_ clknet_leaf_66_wb_clk_i as2650.r0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6648__A2 _1855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6263_ _1630_ _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8002_ _1467_ _3231_ _3233_ _3236_ _3237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_5214_ _0562_ _0567_ _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6194_ _1558_ _1566_ _1570_ _0069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_135_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5145_ _0550_ _0581_ _0584_ _0447_ _0585_ _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_96_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8270__B2 _3472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5076_ _0517_ _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5959__I _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8335__I _3505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8904_ _0065_ clknet_leaf_61_wb_clk_i as2650.r123_2\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_65_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8022__A1 _4322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8835_ _3996_ _3998_ _3049_ _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_77_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_50_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8573__A2 _3765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5387__A2 _4417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6584__A1 _4061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8766_ _1713_ _1048_ _3938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5978_ _1268_ _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7717_ _2824_ _2931_ _2962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4929_ _4375_ _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5694__I _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8697_ _2354_ _1227_ _1245_ _2314_ _3871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__9166__I net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8070__I _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5139__A2 _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6336__A1 _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7648_ _2687_ _2894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7579_ _2777_ _2792_ _2826_ _2732_ _2827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_88_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8089__A1 _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6639__A2 _1960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7064__A2 _2343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4822__A1 _4393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6575__A1 _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6327__A1 _1629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6878__A2 _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7827__A1 _3051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5302__A2 _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5853__A3 _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7260__S _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7055__A2 _2336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5066__A1 _4179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6950_ _1021_ _2218_ _2244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8004__A1 _4079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5901_ _1213_ _1277_ _1292_ _1295_ _0051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_35_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6881_ _1800_ _2187_ _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_78_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8555__A2 _3725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8620_ _2898_ _3807_ _3812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5832_ _4079_ _1226_ _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_8551_ _3089_ _3740_ _3746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5763_ _1143_ _1164_ _1172_ _0036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8307__A2 _4271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7502_ as2650.addr_buff\[1\] _2415_ _2751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4714_ _4115_ _4295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_8482_ _3672_ _3679_ _3579_ _3680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7515__B1 _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5694_ _1120_ _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7515__C2 _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7433_ _2424_ _2663_ _2666_ _2682_ _2683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_136_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4645_ _4225_ _4197_ _4226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5019__I _4302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7364_ _2559_ _2620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4576_ as2650.holding_reg\[0\] _4153_ _4154_ _4157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9103_ _0264_ clknet_leaf_13_wb_clk_i net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7818__A1 _2781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6315_ _1661_ _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7295_ _1237_ _2549_ _1230_ _2554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9034_ _0195_ clknet_leaf_41_wb_clk_i as2650.psu\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__8491__A1 _3667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7294__A2 _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6246_ _1606_ _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6177_ _0784_ _1553_ _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_97_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7046__A2 _2315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5128_ _0468_ _0568_ _0569_ _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_57_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8992__CLK clknet_leaf_46_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5059_ _0490_ _0426_ _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_85_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8818_ _2515_ _3982_ _3984_ _4206_ _3985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_52_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7754__B1 _2691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6021__A3 _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8749_ _2299_ _3920_ _3921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_139_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6309__A1 _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5780__A2 _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7853__B _3093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5532__A2 _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7144__I _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7285__A2 _2539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_36_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_36_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_122_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_110_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8785__A2 _3952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5599__A2 _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6796__A1 _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5220__A1 _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4654__S0 as2650.ins_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6223__I _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8578__C _2629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4430_ _4010_ _4011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__8865__CLK clknet_leaf_58_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5523__A2 _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7054__I _2335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6100_ _0910_ _1403_ _1484_ _1485_ _1486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_112_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8473__A1 _3667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7080_ _2359_ _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7276__A2 _2534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8594__B _3506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5287__A1 _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6031_ _1417_ _1341_ _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6787__A1 _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7982_ _1034_ _2690_ _3208_ _2689_ _3217_ _3218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_81_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7938__B _3175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6933_ _1978_ _2229_ _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_70_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_78_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8528__A2 _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8613__I net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6539__A1 _1855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6864_ _1632_ _2169_ _2171_ as2650.stack\[0\]\[3\] _2174_ _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_126_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8603_ _3790_ _3793_ _3795_ _3602_ _2458_ _3796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__7200__A2 _4292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5815_ _1142_ _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6003__A3 _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6795_ _2081_ _2086_ _2112_ _2113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5211__A1 _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6133__I _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8534_ _0783_ _0796_ _3730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5746_ _1161_ _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5762__A2 _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8465_ _3040_ _2975_ _3493_ _3662_ _3663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5972__I _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5677_ as2650.pc\[9\] _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_136_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7503__A3 _2751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8700__A2 _1846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7416_ _2345_ _2664_ _2665_ _0876_ _2666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_4628_ _4208_ _4209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8396_ _2405_ _3596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5514__A2 _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5193__B _4179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4588__I _4157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7347_ _1438_ _1230_ _2603_ _2604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_104_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4559_ _4065_ _4140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8464__A1 _2804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7267__A2 _2517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7278_ _2430_ _2536_ _2537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_131_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_9017_ _0178_ clknet_leaf_7_wb_clk_i as2650.holding_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6229_ _1067_ _1068_ _1071_ _1080_ _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_89_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8216__A1 _1646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8767__A2 _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6308__I _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5450__A1 _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5202__A1 _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5753__A2 _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6950__A1 _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5505__A2 _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6702__A1 _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7258__A2 _2489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8207__A1 _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8758__A2 _3282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6218__I _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5122__I as2650.r0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6769__A1 _1937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7966__B1 _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7430__A2 _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7718__B1 _2960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5600_ _1031_ _1032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_108_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6580_ _1869_ _1873_ _1902_ _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor3_1
XFILLER_125_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6941__A1 as2650.r123_2\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5744__A2 _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5531_ _0909_ _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8250_ _2284_ _2266_ _1562_ _3454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7497__A2 _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5462_ _0899_ _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7201_ _2471_ _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__9043__CLK clknet_leaf_29_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8181_ as2650.stack\[6\]\[5\] _3393_ _3403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5393_ _0760_ _0831_ _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_7132_ _2269_ _2403_ _2404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7063_ _2343_ _2344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6014_ _1400_ _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5680__A1 _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8749__A2 _3920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5680__B2 as2650.r123_2\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5967__I _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7965_ _3195_ _3201_ _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6916_ _0925_ _2212_ _2214_ _2215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4786__A3 _4365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7896_ _2779_ _3133_ _2770_ _3136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_63_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7185__A1 net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6847_ _1964_ _2162_ _2163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5735__A2 _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6778_ _0649_ _2096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8517_ _2338_ _3714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5729_ as2650.stack\[5\]\[8\] _1151_ _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_143_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7488__A2 _2736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8448_ _3571_ _3646_ _3647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8379_ _3570_ _3578_ _3579_ _3580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5651__B _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6999__A1 _2285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7660__A2 _2903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7412__A2 _2535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5877__I _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4781__I _4088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7176__A1 _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_70_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9066__CLK clknet_leaf_42_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_51_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_51_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__8676__A1 _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7479__A2 _2688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5561__B _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4956__I _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7332__I _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7100__A1 _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5662__A1 _4129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_37_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8600__A1 _3596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7403__A2 _2611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4691__I _4271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6462__I0 _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8163__I _3389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7750_ _2857_ _2985_ _2993_ _2592_ _2994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4962_ _4142_ _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6701_ _0452_ _1966_ _1907_ _2020_ _2021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_7681_ _2338_ _2927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4893_ _0336_ _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6632_ _1948_ _1953_ _1954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_137_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6563_ _0592_ _0369_ _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8112__B _2547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8302_ _2269_ _2270_ _2271_ _3505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_118_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5514_ as2650.stack\[3\]\[9\] _0948_ _0950_ _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6411__I _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8667__A1 _3838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6494_ _4202_ _1813_ _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8233_ as2650.stack\[7\]\[10\] _3440_ _3442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5445_ _4109_ _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5027__I _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8419__A1 _2910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8164_ _1598_ _3388_ _3390_ as2650.stack\[6\]\[0\] _3385_ _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__7890__A2 _3125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5376_ _0410_ _0801_ _0813_ _0814_ _4147_ _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_4
XFILLER_114_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7115_ _4250_ _2387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_82_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8095_ _2261_ _3326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7046_ _2314_ _2315_ _2328_ _2254_ _2329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_102_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5653__A1 _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8997_ _0158_ clknet_leaf_11_wb_clk_i as2650.addr_buff\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5405__A1 as2650.r0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7948_ _3029_ _3185_ _2465_ _3186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_103_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9089__CLK clknet_leaf_26_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7879_ _3118_ _3119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_51_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6905__A1 _2163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5708__A2 _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__8658__A1 _3838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7330__A1 _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8926__CLK clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7330__B2 _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7094__B1 _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7633__A2 _2877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4447__A2 as2650.cycle\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6991__I _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8189__A3 _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7397__A1 _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7149__A1 _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6231__I _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8649__A1 _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6124__A2 _4241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5230_ _0336_ _0368_ _0466_ _4381_ _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_142_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5291__B _4258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5161_ _0601_ _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7062__I _2276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7085__B1 _2364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8821__A1 _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5092_ _0533_ _4021_ _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6832__B1 _2147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8920_ _0081_ clknet_leaf_32_wb_clk_i as2650.stack\[5\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_42_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8851_ _0012_ clknet_leaf_66_wb_clk_i as2650.r123\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_25_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8585__B1 _3493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8107__B _3337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_40_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7802_ _2832_ _3011_ _3019_ _2842_ _3044_ _3045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__6406__I _1744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5994_ _1365_ _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8782_ _3951_ _1261_ _3953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6060__A1 _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4945_ _0387_ _0294_ _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7733_ _2882_ _2976_ _2894_ _2977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_127_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7664_ _1410_ _2809_ _2910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4876_ _0319_ _4388_ _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_71_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6899__B1 _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6615_ _0588_ _1936_ _1937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7595_ _2690_ _2842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8949__CLK clknet_leaf_34_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6363__A2 _1592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7237__I _2490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6141__I _4078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6546_ _0820_ _0856_ _1868_ _1869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_10_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5571__B1 _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7312__A1 _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6477_ _1797_ _4314_ _1799_ _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__6115__A2 _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5428_ _4111_ _0864_ _0865_ _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_8216_ _1646_ _3416_ _3417_ _3430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5874__A1 _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5359_ _4368_ _0797_ _0293_ _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_8147_ _0887_ _3019_ _3374_ _3282_ _3375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8078_ _3277_ _0458_ _3310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8812__A1 _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7029_ _2312_ _1586_ _2294_ _2313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7379__A1 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8040__A2 _4186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5929__A2 _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output14_I net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4601__A2 _4156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7551__A1 _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7303__A1 _2311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5890__I _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__9104__CLK clknet_leaf_13_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7606__A2 _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6409__A3 _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8803__A1 _1475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7610__I _2704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4840__A2 _4322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8031__A2 _4250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4979__I0 as2650.r123\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7790__A1 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4730_ _4310_ _4192_ _4311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4661_ _4241_ _4242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7542__A1 _2782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7057__I _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7542__B2 _2788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6400_ _1649_ _1712_ _1740_ _0105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7380_ _2633_ _2634_ _2339_ _2635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_70_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4592_ as2650.carry _4173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__8597__B _3472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6331_ _1689_ _1672_ _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_128_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8098__A2 _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_7_wb_clk_i_I clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_9050_ _0211_ clknet_leaf_64_wb_clk_i as2650.r0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6262_ as2650.pc\[3\] _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8001_ _1420_ _3235_ _3236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5213_ _0576_ _0653_ _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6193_ _1569_ _1563_ _1555_ _1549_ _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_130_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5144_ _4270_ _0535_ _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6845__B _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5075_ _0418_ _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6281__A1 _1646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8903_ _0064_ clknet_leaf_73_wb_clk_i as2650.r123_2\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6281__B2 as2650.stack\[5\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8022__A2 _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8834_ _2519_ _3997_ _3998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6033__A1 _4292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8573__A3 _3766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8765_ _2603_ _3937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5975__I _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5387__A3 _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6584__A2 _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5977_ _4224_ _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_80_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4595__A1 _4175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7716_ _2823_ _2961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4928_ _4415_ _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8696_ _3869_ _1576_ _3870_ _0271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7647_ _2885_ _2881_ _2890_ _2892_ _2758_ _2893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_100_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7533__A1 _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4859_ _4190_ _0301_ _0302_ _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__5139__A3 _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7578_ _2790_ _2815_ _2822_ _2823_ _2825_ _2826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_119_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6529_ _1851_ _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8089__A2 _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7836__A2 _3053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6046__I _4084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7772__A1 _3012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8261__I _4365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4586__A1 _4166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6327__A2 _1662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7524__A1 _1615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4510__A1 _4090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7055__A3 _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8004__A2 _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5900_ _1294_ _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6880_ _1542_ _1862_ _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_62_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5831_ _1223_ _1225_ _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5795__I _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7763__A1 _2968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7763__B2 _2688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4577__A1 _4156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8550_ _3625_ _3744_ _3745_ _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5762_ as2650.stack\[6\]\[14\] _1162_ _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8104__C _2586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7501_ _4393_ _1072_ _2750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4713_ _4293_ _4294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8481_ _3603_ _3677_ _3678_ _2287_ _3679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5693_ as2650.pc\[11\] _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7515__B2 as2650.stack\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7432_ _2671_ _2674_ _2679_ _2681_ _2682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_15_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4644_ _4080_ _4072_ _4225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_129_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7363_ _2542_ _1071_ _2617_ _2618_ _2619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4575_ _4113_ _4153_ _4155_ _4156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_116_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8120__B _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_9102_ _0263_ clknet_leaf_13_wb_clk_i net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6314_ _1619_ _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7294_ _2547_ _2319_ _2549_ _2552_ _2553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__7818__A2 _3053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9033_ _0194_ clknet_leaf_17_wb_clk_i as2650.cycle\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6245_ _1614_ _1615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_103_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4501__A1 _4034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6176_ _4105_ _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_83_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5127_ _0417_ _4319_ _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5058_ _0495_ _0498_ _0499_ _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_38_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8817_ _2303_ _2517_ _3978_ _3984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7754__A1 as2650.stack\[7\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8081__I _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8748_ _2421_ _3920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6021__A4 _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8679_ _3851_ _3857_ _3858_ _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7506__A1 _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6309__A2 _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7853__C _2789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5373__C _4348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_49_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7285__A3 _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5296__A2 _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8256__I _3459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8234__A2 _3437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_76_wb_clk_i clknet_3_0_0_wb_clk_i clknet_leaf_76_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_114_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7993__A1 _2652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6796__A2 _2076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4654__S1 _4010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7335__I _2464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4731__A1 _4297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6484__A1 _4366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6030_ _4040_ _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input5_I io_in[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7981_ _2461_ _3215_ _3216_ _3217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_67_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7984__A1 as2650.pc\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6932_ _2207_ _2229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7938__C _2758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_63_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4643__B _4175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6863_ _1620_ _2167_ _2175_ _0133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7736__A1 _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6539__A2 _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8602_ _3147_ _3794_ _3795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_23_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5814_ _1209_ _1198_ _1210_ _0049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6794_ _0588_ _2076_ _2087_ _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_37_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_8533_ _2252_ _3728_ _3729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7954__B _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5745_ _1145_ _1160_ _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_124_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8464_ _2804_ _3661_ _2980_ _3662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5676_ _1087_ _1103_ _1105_ _0016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_135_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7415_ _1463_ _2276_ _2665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4627_ as2650.r0\[7\] _4208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8395_ _2532_ _3595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4722__A1 _4285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7346_ _1273_ _2603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_11_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4558_ _4135_ _4139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_117_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8785__B _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8464__A2 _3661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7277_ _1546_ _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4489_ _4069_ _4070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_104_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6475__A1 _4286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5278__A2 _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_9016_ _0177_ clknet_leaf_10_wb_clk_i as2650.idx_ctrl\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6228_ _1598_ _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6159_ as2650.r123_2\[3\]\[5\] _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__9112__D _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7975__A1 as2650.pc\[14\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7727__A1 as2650.pc\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5202__A2 _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4961__A1 _4343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4961__B2 _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8152__A1 _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7155__I _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput40 net40 io_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_64_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6466__A1 _1738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7966__A1 _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7966__B2 _2996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7430__A3 _2265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7718__B2 _2961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6234__I _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8391__A1 _3581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5530_ _4017_ _0965_ _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__8143__A1 _3340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5461_ _0898_ _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7497__A3 _2734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7200_ _1242_ _4292_ _2471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5392_ as2650.r0\[6\] _4414_ _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8180_ _2177_ _3398_ _3401_ _3402_ _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_114_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7131_ _4090_ _2270_ _2271_ _2403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_125_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6457__A1 _1629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7062_ _2276_ _2343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6013_ _4392_ _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6209__A1 _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6209__B2 _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7957__A1 _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7421__A3 _2667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7964_ _2857_ _3197_ _3194_ _2882_ _3200_ _3201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6915_ _0876_ _1799_ _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7709__A1 _2857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7895_ _0980_ _2842_ _3113_ _2832_ _3134_ _3135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_6846_ _2159_ _2160_ _2161_ _2162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7185__A2 _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5196__A1 _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6777_ _1962_ _2068_ _2070_ _2095_ _0127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5983__I _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8516_ _3459_ _3713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5728_ _1149_ _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4943__A1 _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__8134__A1 _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_8447_ _3640_ _3641_ _3644_ _3646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_87_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5659_ _1051_ _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8685__A2 _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6696__A1 _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8378_ _2404_ _3579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7329_ _2584_ _2585_ _2586_ _2587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_132_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6999__A2 _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5120__A1 _4148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6319__I _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7660__A3 _2904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7859__B _4293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7948__A1 _3029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6620__A1 as2650.r0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8855__CLK clknet_leaf_47_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8373__A1 _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7176__A2 _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6989__I _4293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4934__A1 _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8125__A1 _3339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7613__I _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6439__A1 as2650.stack\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5662__A2 _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7939__A1 _2882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4972__I _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_30_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6462__I1 as2650.stack\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4961_ _4343_ _0394_ _0402_ _0403_ _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_45_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6700_ _2018_ _2019_ _1918_ _2020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_75_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7680_ _2881_ _2895_ _2925_ _2688_ _2926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_75_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4892_ _0335_ _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6631_ _1950_ _1952_ _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_60_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6562_ _0841_ _0851_ _1884_ _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8116__A1 as2650.psl\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8301_ _1400_ _3465_ _3504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5513_ _0949_ _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__8667__A2 _2014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6127__B1 _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6493_ _1815_ _1816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8232_ _1200_ _3437_ _3441_ _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_121_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5444_ _0881_ _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5350__A1 _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8163_ _3389_ _3390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5375_ _0405_ _0800_ _4164_ _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_99_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7627__B1 _2841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7114_ _4088_ _4027_ _4400_ _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_87_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8094_ _3271_ _0516_ _3324_ _3325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7045_ _1062_ _1431_ _2317_ _2327_ _2328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_68_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8878__CLK clknet_leaf_58_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6850__A1 _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5653__A2 _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8996_ _0157_ clknet_leaf_23_wb_clk_i as2650.addr_buff\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_23_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7947_ _1129_ _3184_ _3185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_97_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8355__A1 _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7878_ as2650.pc\[10\] _2987_ _3118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_51_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8355__B2 _3294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5169__A1 _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6829_ _0701_ _1848_ _2145_ _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6905__A2 _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4916__A1 _4252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8107__A1 _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6118__B1 _4389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8658__A2 _3262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6669__A1 _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4931__A4 _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5341__A1 _4222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5341__B2 _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5154__S _4013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7094__A1 _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6841__A1 _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5888__I _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6444__I1 _4306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__9033__CLK clknet_leaf_17_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8346__A1 _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7149__A2 _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4907__A1 _4063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8649__A2 _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4967__I _4331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5160_ _0600_ _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_123_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7085__A1 _4317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8282__B1 _3484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5091_ as2650.r0\[5\] _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5635__A2 _4124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6832__A1 _2013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6832__B2 _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8850_ _0011_ clknet_leaf_67_wb_clk_i as2650.r123\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7388__A2 _2637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8585__A1 _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8107__C _2730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8585__B2 _3778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7801_ _3028_ _3041_ _3042_ _3043_ _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_65_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5399__A1 as2650.r0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8781_ _1355_ _2657_ _3952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5993_ _0711_ _1260_ _1379_ _0938_ _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_91_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6060__A2 _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7732_ _2885_ _2968_ _2975_ _2892_ _2758_ _2976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_4944_ as2650.holding_reg\[2\] _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__8337__A1 _4392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_33_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7663_ _2793_ _2908_ _2909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__8123__B _3352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4875_ _4160_ _4232_ _4234_ _4236_ _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__6899__A1 _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6614_ _1935_ _1936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7594_ _2840_ _2841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_118_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7962__B _3198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6545_ _0825_ _0855_ _1868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6476_ _1798_ _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7312__A2 _2535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8215_ as2650.stack\[7\]\[5\] _3413_ _3429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5427_ _4093_ _4091_ _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5323__A1 as2650.r0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7253__I _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8146_ _1518_ _3283_ _3373_ _3374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5358_ _0796_ _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7076__A1 _2347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8077_ _3271_ _0452_ _3309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5289_ _4380_ _0714_ _0728_ _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5626__A2 _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6823__A1 _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7028_ _2311_ _2312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_74_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__9056__CLK clknet_leaf_67_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8025__B1 _4224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__8576__A1 net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7379__A2 _2613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8979_ _0140_ clknet_leaf_3_wb_clk_i as2650.r123_2\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_83_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6051__A2 _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__8328__A1 _2884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7000__A1 _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5376__C _4147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7551__A2 _2593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7303__A2 _2561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8500__A1 _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8259__I _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5314__A1 _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7067__A1 _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8803__A2 _3906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7112__B _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6042__A2 _4125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4979__I1 as2650.r123\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8319__A1 _1615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__8319__B2 _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7790__A2 _4215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5567__B _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6242__I as2650.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4660_ net5 _4241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7542__A2 _2777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4591_ _4141_ _4171_ _4172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6330_ _1688_ _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_127_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5305__A1 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5156__I1 as2650.r123\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6261_ _1628_ _1629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_89_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7073__I _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8000_ _1078_ _3234_ _3235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5212_ _0559_ _0574_ _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6192_ _1568_ _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7058__A1 net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5143_ _0582_ _0583_ _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_9_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5074_ _0515_ _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_8902_ _0063_ clknet_leaf_71_wb_clk_i as2650.r123_2\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_38_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8833_ _3952_ _3991_ _3997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6569__B1 _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7230__A1 _4194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6033__A2 _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8916__CLK clknet_leaf_33_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8764_ _3921_ _3935_ _3936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5976_ _4101_ _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7715_ _2955_ _2957_ _2958_ _2959_ _2960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_4927_ _4187_ _0370_ _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_8695_ _2307_ _1573_ _3870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7248__I _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7646_ _2891_ _2892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4858_ as2650.holding_reg\[2\] _4190_ _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7533__A2 _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5139__A4 _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7692__B _2936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7577_ _2824_ _2777_ _2825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4789_ _4257_ _4369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6528_ _1520_ _1850_ _1851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_109_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7297__A1 _2537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7297__B2 _2431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6459_ _1689_ _1782_ _1785_ _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_122_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7049__A1 _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_8129_ _3340_ _0735_ _2898_ _3358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7711__I _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7772__A2 _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5783__A1 _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4586__A2 _4143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7158__I _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6062__I _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7524__A2 _2731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8210__C _3409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8485__B1 _3682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5838__A2 _4004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4510__A2 _4055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7621__I _2809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7055__A4 _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7460__A1 _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8939__CLK clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6237__I _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5830_ _1224_ _4128_ _4145_ _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_61_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5761_ _1138_ _1164_ _1171_ _0035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_61_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4577__A2 _4157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7500_ _2711_ _2748_ _2749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4712_ _4292_ _4293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_8480_ _0726_ _3544_ _3678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5692_ _1087_ _1118_ _1119_ _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__8712__A1 _3313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7431_ _2401_ _2452_ _2618_ _2680_ _2681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_124_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5526__A1 _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4643_ _4207_ _4223_ _4175_ _4224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_102_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7362_ _0784_ _2353_ _1545_ _2618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_128_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4574_ as2650.holding_reg\[0\] _4154_ _4155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_144_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_9101_ _0262_ clknet_leaf_13_wb_clk_i net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7279__A1 _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6313_ _1611_ _1662_ _1674_ _0084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7293_ _1560_ _2550_ _2551_ _1229_ _2552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_9032_ _0193_ clknet_leaf_23_wb_clk_i as2650.cycle\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6244_ _1613_ _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4501__A2 _4081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6175_ _1427_ _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_69_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__8779__A1 _3935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5126_ _0336_ _4415_ _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_69_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5057_ _0495_ _0498_ _0385_ _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5986__I _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7203__A1 _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4890__I _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8816_ _2533_ _3983_ _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8747_ _3910_ _3918_ _3919_ _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_90_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5959_ _1345_ _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_80_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_8678_ net45 _3846_ _3858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7506__A2 _2749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8703__A1 _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5935__B _4344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7629_ _2834_ _2875_ _2876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_5_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7441__I _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7993__A2 _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_45_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_72_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6520__I _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6181__A1 _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4731__A2 _4300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4975__I _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6484__A2 _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_141_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_39_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7980_ _2701_ _2778_ _3208_ _3216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__9117__CLK clknet_leaf_66_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7984__A2 _2731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6931_ as2650.r123_2\[0\]\[2\] _2224_ _2227_ _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5995__A1 _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6862_ _1624_ _2169_ _2171_ as2650.stack\[0\]\[2\] _2174_ _2175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_81_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7736__A2 _2851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8601_ _3120_ _3774_ _3148_ _3794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_39_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5813_ as2650.stack\[1\]\[13\] _1196_ _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6793_ _2109_ _2093_ _2110_ _2111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_8532_ _3725_ _3727_ _3728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5744_ _1146_ _0908_ _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_8463_ net34 _3660_ _3661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5675_ as2650.stack\[3\]\[8\] _1104_ _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7414_ _1858_ _2355_ _2664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4626_ _4206_ _4207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_8394_ _3489_ _3593_ _3594_ _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7345_ _1055_ _2592_ _2597_ _2601_ _2602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_116_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4557_ _4137_ _4138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4722__A2 _4302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7276_ _2334_ _2534_ _2535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4488_ as2650.ins_reg\[7\] _4069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_9015_ _0176_ clknet_leaf_10_wb_clk_i as2650.idx_ctrl\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6475__A2 _4110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5278__A3 _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6227_ _1597_ _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6158_ _1538_ _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_100_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7424__A1 _4362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5109_ _0443_ _0425_ _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_46_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6089_ _0804_ _0815_ _1475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_3427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7975__A2 _3210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7727__A2 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__8025__C _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_41_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7864__C _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7436__I _2685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput30 net30 io_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput41 net41 io_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_107_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7663__A1 _2793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4795__I _4229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6466__A2 _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7415__A1 _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_97_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7966__A2 _2961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8143__A2 _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7346__I _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6250__I _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5460_ _0895_ _0897_ _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_121_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5391_ _0668_ _0672_ _0829_ _0821_ _0755_ _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_1
XFILLER_119_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7130_ _2400_ _2401_ _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__8446__A3 _3644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7654__A1 _2899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6457__A2 _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7061_ _2275_ _2341_ _2342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7081__I _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6012_ _1398_ _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
.ends

