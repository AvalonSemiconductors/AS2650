magic
tech gf180mcuD
magscale 1 5
timestamp 1701963768
<< obsm1 >>
rect 672 1538 20328 19305
<< metal2 >>
rect 1232 20600 1288 21000
rect 2912 20600 2968 21000
rect 4592 20600 4648 21000
rect 6272 20600 6328 21000
rect 7952 20600 8008 21000
rect 9632 20600 9688 21000
rect 11312 20600 11368 21000
rect 12992 20600 13048 21000
rect 14672 20600 14728 21000
rect 16352 20600 16408 21000
rect 18032 20600 18088 21000
rect 19712 20600 19768 21000
<< obsm2 >>
rect 574 20570 1202 20650
rect 1318 20570 2882 20650
rect 2998 20570 4562 20650
rect 4678 20570 6242 20650
rect 6358 20570 7922 20650
rect 8038 20570 9602 20650
rect 9718 20570 11282 20650
rect 11398 20570 12962 20650
rect 13078 20570 14642 20650
rect 14758 20570 16322 20650
rect 16438 20570 18002 20650
rect 18118 20570 19682 20650
rect 574 1549 19754 20570
<< metal3 >>
rect 0 19152 400 19208
rect 0 18704 400 18760
rect 0 18256 400 18312
rect 0 17808 400 17864
rect 0 17360 400 17416
rect 0 16912 400 16968
rect 0 16464 400 16520
rect 0 16016 400 16072
rect 0 15568 400 15624
rect 0 15120 400 15176
rect 0 14672 400 14728
rect 0 14224 400 14280
rect 0 13776 400 13832
rect 0 13328 400 13384
rect 0 12880 400 12936
rect 0 12432 400 12488
rect 0 11984 400 12040
rect 0 11536 400 11592
rect 0 11088 400 11144
rect 0 10640 400 10696
rect 0 10192 400 10248
rect 0 9744 400 9800
rect 0 9296 400 9352
rect 0 8848 400 8904
rect 0 8400 400 8456
rect 0 7952 400 8008
rect 0 7504 400 7560
rect 0 7056 400 7112
rect 0 6608 400 6664
rect 0 6160 400 6216
rect 0 5712 400 5768
rect 0 5264 400 5320
rect 0 4816 400 4872
rect 0 4368 400 4424
rect 0 3920 400 3976
rect 0 3472 400 3528
rect 0 3024 400 3080
rect 0 2576 400 2632
rect 0 2128 400 2184
rect 0 1680 400 1736
<< obsm3 >>
rect 430 19122 18863 19222
rect 400 18790 18863 19122
rect 430 18674 18863 18790
rect 400 18342 18863 18674
rect 430 18226 18863 18342
rect 400 17894 18863 18226
rect 430 17778 18863 17894
rect 400 17446 18863 17778
rect 430 17330 18863 17446
rect 400 16998 18863 17330
rect 430 16882 18863 16998
rect 400 16550 18863 16882
rect 430 16434 18863 16550
rect 400 16102 18863 16434
rect 430 15986 18863 16102
rect 400 15654 18863 15986
rect 430 15538 18863 15654
rect 400 15206 18863 15538
rect 430 15090 18863 15206
rect 400 14758 18863 15090
rect 430 14642 18863 14758
rect 400 14310 18863 14642
rect 430 14194 18863 14310
rect 400 13862 18863 14194
rect 430 13746 18863 13862
rect 400 13414 18863 13746
rect 430 13298 18863 13414
rect 400 12966 18863 13298
rect 430 12850 18863 12966
rect 400 12518 18863 12850
rect 430 12402 18863 12518
rect 400 12070 18863 12402
rect 430 11954 18863 12070
rect 400 11622 18863 11954
rect 430 11506 18863 11622
rect 400 11174 18863 11506
rect 430 11058 18863 11174
rect 400 10726 18863 11058
rect 430 10610 18863 10726
rect 400 10278 18863 10610
rect 430 10162 18863 10278
rect 400 9830 18863 10162
rect 430 9714 18863 9830
rect 400 9382 18863 9714
rect 430 9266 18863 9382
rect 400 8934 18863 9266
rect 430 8818 18863 8934
rect 400 8486 18863 8818
rect 430 8370 18863 8486
rect 400 8038 18863 8370
rect 430 7922 18863 8038
rect 400 7590 18863 7922
rect 430 7474 18863 7590
rect 400 7142 18863 7474
rect 430 7026 18863 7142
rect 400 6694 18863 7026
rect 430 6578 18863 6694
rect 400 6246 18863 6578
rect 430 6130 18863 6246
rect 400 5798 18863 6130
rect 430 5682 18863 5798
rect 400 5350 18863 5682
rect 430 5234 18863 5350
rect 400 4902 18863 5234
rect 430 4786 18863 4902
rect 400 4454 18863 4786
rect 430 4338 18863 4454
rect 400 4006 18863 4338
rect 430 3890 18863 4006
rect 400 3558 18863 3890
rect 430 3442 18863 3558
rect 400 3110 18863 3442
rect 430 2994 18863 3110
rect 400 2662 18863 2994
rect 430 2546 18863 2662
rect 400 2214 18863 2546
rect 430 2098 18863 2214
rect 400 1766 18863 2098
rect 430 1650 18863 1766
rect 400 1554 18863 1650
<< metal4 >>
rect 2224 1538 2384 19238
rect 9904 1538 10064 19238
rect 17584 1538 17744 19238
<< obsm4 >>
rect 1190 4041 2194 18975
rect 2414 4041 9874 18975
rect 10094 4041 12138 18975
<< labels >>
rlabel metal2 s 7952 20600 8008 21000 6 bus_out[0]
port 1 nsew signal output
rlabel metal2 s 9632 20600 9688 21000 6 bus_out[1]
port 2 nsew signal output
rlabel metal2 s 11312 20600 11368 21000 6 bus_out[2]
port 3 nsew signal output
rlabel metal2 s 12992 20600 13048 21000 6 bus_out[3]
port 4 nsew signal output
rlabel metal2 s 14672 20600 14728 21000 6 bus_out[4]
port 5 nsew signal output
rlabel metal2 s 16352 20600 16408 21000 6 bus_out[5]
port 6 nsew signal output
rlabel metal2 s 18032 20600 18088 21000 6 bus_out[6]
port 7 nsew signal output
rlabel metal2 s 19712 20600 19768 21000 6 bus_out[7]
port 8 nsew signal output
rlabel metal2 s 2912 20600 2968 21000 6 cs_port[0]
port 9 nsew signal input
rlabel metal2 s 4592 20600 4648 21000 6 cs_port[1]
port 10 nsew signal input
rlabel metal2 s 6272 20600 6328 21000 6 cs_port[2]
port 11 nsew signal input
rlabel metal3 s 0 16016 400 16072 6 last_addr[0]
port 12 nsew signal input
rlabel metal3 s 0 16464 400 16520 6 last_addr[1]
port 13 nsew signal input
rlabel metal3 s 0 16912 400 16968 6 last_addr[2]
port 14 nsew signal input
rlabel metal3 s 0 17360 400 17416 6 last_addr[3]
port 15 nsew signal input
rlabel metal3 s 0 17808 400 17864 6 last_addr[4]
port 16 nsew signal input
rlabel metal3 s 0 18256 400 18312 6 last_addr[5]
port 17 nsew signal input
rlabel metal3 s 0 18704 400 18760 6 last_addr[6]
port 18 nsew signal input
rlabel metal3 s 0 19152 400 19208 6 last_addr[7]
port 19 nsew signal input
rlabel metal3 s 0 8848 400 8904 6 ram_end[0]
port 20 nsew signal input
rlabel metal3 s 0 13328 400 13384 6 ram_end[10]
port 21 nsew signal input
rlabel metal3 s 0 13776 400 13832 6 ram_end[11]
port 22 nsew signal input
rlabel metal3 s 0 14224 400 14280 6 ram_end[12]
port 23 nsew signal input
rlabel metal3 s 0 14672 400 14728 6 ram_end[13]
port 24 nsew signal input
rlabel metal3 s 0 15120 400 15176 6 ram_end[14]
port 25 nsew signal input
rlabel metal3 s 0 15568 400 15624 6 ram_end[15]
port 26 nsew signal input
rlabel metal3 s 0 9296 400 9352 6 ram_end[1]
port 27 nsew signal input
rlabel metal3 s 0 9744 400 9800 6 ram_end[2]
port 28 nsew signal input
rlabel metal3 s 0 10192 400 10248 6 ram_end[3]
port 29 nsew signal input
rlabel metal3 s 0 10640 400 10696 6 ram_end[4]
port 30 nsew signal input
rlabel metal3 s 0 11088 400 11144 6 ram_end[5]
port 31 nsew signal input
rlabel metal3 s 0 11536 400 11592 6 ram_end[6]
port 32 nsew signal input
rlabel metal3 s 0 11984 400 12040 6 ram_end[7]
port 33 nsew signal input
rlabel metal3 s 0 12432 400 12488 6 ram_end[8]
port 34 nsew signal input
rlabel metal3 s 0 12880 400 12936 6 ram_end[9]
port 35 nsew signal input
rlabel metal3 s 0 1680 400 1736 6 ram_start[0]
port 36 nsew signal input
rlabel metal3 s 0 6160 400 6216 6 ram_start[10]
port 37 nsew signal input
rlabel metal3 s 0 6608 400 6664 6 ram_start[11]
port 38 nsew signal input
rlabel metal3 s 0 7056 400 7112 6 ram_start[12]
port 39 nsew signal input
rlabel metal3 s 0 7504 400 7560 6 ram_start[13]
port 40 nsew signal input
rlabel metal3 s 0 7952 400 8008 6 ram_start[14]
port 41 nsew signal input
rlabel metal3 s 0 8400 400 8456 6 ram_start[15]
port 42 nsew signal input
rlabel metal3 s 0 2128 400 2184 6 ram_start[1]
port 43 nsew signal input
rlabel metal3 s 0 2576 400 2632 6 ram_start[2]
port 44 nsew signal input
rlabel metal3 s 0 3024 400 3080 6 ram_start[3]
port 45 nsew signal input
rlabel metal3 s 0 3472 400 3528 6 ram_start[4]
port 46 nsew signal input
rlabel metal3 s 0 3920 400 3976 6 ram_start[5]
port 47 nsew signal input
rlabel metal3 s 0 4368 400 4424 6 ram_start[6]
port 48 nsew signal input
rlabel metal3 s 0 4816 400 4872 6 ram_start[7]
port 49 nsew signal input
rlabel metal3 s 0 5264 400 5320 6 ram_start[8]
port 50 nsew signal input
rlabel metal3 s 0 5712 400 5768 6 ram_start[9]
port 51 nsew signal input
rlabel metal4 s 2224 1538 2384 19238 6 vdd
port 52 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 19238 6 vdd
port 52 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 19238 6 vss
port 53 nsew ground bidirectional
rlabel metal2 s 1232 20600 1288 21000 6 wb_clk_i
port 54 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 21000 21000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1140074
string GDS_FILE /run/media/tholin/fbc90f8f-67e9-406d-9872-54f02ad6a2d8/AS2650/openlane/boot_rom/runs/23_12_07_16_40/results/signoff/boot_rom.magic.gds
string GDS_START 295462
<< end >>

