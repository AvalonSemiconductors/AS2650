VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO avali_logo
  CLASS BLOCK ;
  FOREIGN avali_logo ;
  ORIGIN 0.000 0.000 ;
  SIZE 375.000 BY 440.250 ;
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal4 ;
        RECT 141.000 302.250 161.250 303.000 ;
        RECT 133.500 301.500 171.000 302.250 ;
        RECT 127.500 300.750 178.500 301.500 ;
        RECT 123.750 300.000 183.750 300.750 ;
        RECT 120.000 299.250 183.750 300.000 ;
        RECT 116.250 298.500 183.000 299.250 ;
        RECT 113.250 297.750 183.000 298.500 ;
        RECT 111.000 297.000 182.250 297.750 ;
        RECT 108.000 296.250 182.250 297.000 ;
        RECT 105.750 295.500 181.500 296.250 ;
        RECT 103.500 294.750 181.500 295.500 ;
        RECT 101.250 294.000 180.750 294.750 ;
        RECT 99.000 293.250 180.000 294.000 ;
        RECT 97.500 292.500 180.000 293.250 ;
        RECT 95.250 291.750 179.250 292.500 ;
        RECT 93.750 291.000 179.250 291.750 ;
        RECT 91.500 290.250 178.500 291.000 ;
        RECT 90.000 289.500 178.500 290.250 ;
        RECT 88.500 288.750 177.750 289.500 ;
        RECT 87.000 288.000 177.750 288.750 ;
        RECT 85.500 287.250 177.000 288.000 ;
        RECT 84.000 286.500 177.000 287.250 ;
        RECT 82.500 285.750 176.250 286.500 ;
        RECT 81.000 285.000 176.250 285.750 ;
        RECT 79.500 284.250 175.500 285.000 ;
        RECT 78.000 283.500 174.750 284.250 ;
        RECT 76.500 282.750 174.750 283.500 ;
        RECT 75.000 282.000 174.000 282.750 ;
        RECT 74.250 281.250 174.000 282.000 ;
        RECT 72.750 280.500 173.250 281.250 ;
        RECT 72.000 279.750 173.250 280.500 ;
        RECT 70.500 279.000 172.500 279.750 ;
        RECT 69.000 278.250 172.500 279.000 ;
        RECT 68.250 277.500 171.750 278.250 ;
        RECT 66.750 276.750 171.750 277.500 ;
        RECT 66.000 276.000 139.500 276.750 ;
        RECT 165.750 276.000 171.000 276.750 ;
        RECT 64.500 275.250 133.500 276.000 ;
        RECT 63.750 274.500 129.000 275.250 ;
        RECT 63.000 273.750 125.250 274.500 ;
        RECT 61.500 273.000 122.250 273.750 ;
        RECT 60.750 272.250 119.250 273.000 ;
        RECT 60.000 271.500 116.250 272.250 ;
        RECT 58.500 270.750 114.000 271.500 ;
        RECT 57.750 270.000 111.750 270.750 ;
        RECT 57.000 269.250 109.500 270.000 ;
        RECT 55.500 268.500 107.250 269.250 ;
        RECT 54.750 267.750 105.750 268.500 ;
        RECT 54.000 267.000 103.500 267.750 ;
        RECT 53.250 266.250 102.000 267.000 ;
        RECT 52.500 265.500 100.500 266.250 ;
        RECT 51.750 264.750 98.250 265.500 ;
        RECT 50.250 264.000 96.750 264.750 ;
        RECT 49.500 263.250 95.250 264.000 ;
        RECT 48.750 262.500 93.750 263.250 ;
        RECT 48.000 261.750 92.250 262.500 ;
        RECT 47.250 261.000 91.500 261.750 ;
        RECT 46.500 260.250 90.000 261.000 ;
        RECT 45.750 259.500 88.500 260.250 ;
        RECT 45.000 258.750 87.000 259.500 ;
        RECT 44.250 258.000 86.250 258.750 ;
        RECT 43.500 257.250 84.750 258.000 ;
        RECT 42.750 256.500 84.000 257.250 ;
        RECT 42.000 255.750 82.500 256.500 ;
        RECT 41.250 255.000 81.000 255.750 ;
        RECT 40.500 254.250 80.250 255.000 ;
        RECT 39.750 253.500 79.500 254.250 ;
        RECT 39.000 252.750 78.000 253.500 ;
        RECT 39.000 252.000 77.250 252.750 ;
        RECT 38.250 251.250 75.750 252.000 ;
        RECT 37.500 250.500 75.000 251.250 ;
        RECT 36.750 249.750 74.250 250.500 ;
        RECT 36.000 249.000 73.500 249.750 ;
        RECT 35.250 248.250 72.000 249.000 ;
        RECT 34.500 247.500 71.250 248.250 ;
        RECT 34.500 246.750 70.500 247.500 ;
        RECT 33.750 246.000 69.750 246.750 ;
        RECT 33.000 245.250 69.000 246.000 ;
        RECT 32.250 244.500 68.250 245.250 ;
        RECT 31.500 243.750 66.750 244.500 ;
        RECT 31.500 243.000 66.000 243.750 ;
        RECT 30.750 242.250 65.250 243.000 ;
        RECT 30.000 241.500 64.500 242.250 ;
        RECT 29.250 240.750 63.750 241.500 ;
        RECT 29.250 240.000 63.000 240.750 ;
        RECT 28.500 239.250 62.250 240.000 ;
        RECT 27.750 238.500 61.500 239.250 ;
        RECT 27.750 237.750 60.750 238.500 ;
        RECT 27.000 237.000 60.000 237.750 ;
        RECT 26.250 236.250 59.250 237.000 ;
        RECT 25.500 234.750 58.500 236.250 ;
        RECT 24.750 234.000 57.750 234.750 ;
        RECT 24.750 233.250 57.000 234.000 ;
        RECT 24.000 232.500 56.250 233.250 ;
        RECT 23.250 231.750 55.500 232.500 ;
        RECT 23.250 231.000 54.750 231.750 ;
        RECT 22.500 230.250 54.000 231.000 ;
        RECT 21.750 229.500 54.000 230.250 ;
        RECT 21.750 228.750 53.250 229.500 ;
        RECT 21.000 228.000 52.500 228.750 ;
        RECT 21.000 227.250 51.750 228.000 ;
        RECT 20.250 226.500 51.750 227.250 ;
        RECT 19.500 225.750 51.000 226.500 ;
        RECT 19.500 225.000 50.250 225.750 ;
        RECT 18.750 223.500 49.500 225.000 ;
        RECT 18.000 222.750 48.750 223.500 ;
        RECT 18.000 222.000 48.000 222.750 ;
        RECT 17.250 221.250 48.000 222.000 ;
        RECT 17.250 220.500 47.250 221.250 ;
        RECT 16.500 219.000 46.500 220.500 ;
        RECT 15.750 218.250 45.750 219.000 ;
        RECT 15.750 217.500 45.000 218.250 ;
        RECT 15.000 216.750 45.000 217.500 ;
        RECT 15.000 216.000 44.250 216.750 ;
        RECT 14.250 214.500 43.500 216.000 ;
        RECT 13.500 213.000 42.750 214.500 ;
        RECT 12.750 211.500 42.000 213.000 ;
        RECT 12.750 210.750 41.250 211.500 ;
        RECT 12.000 210.000 41.250 210.750 ;
        RECT 12.000 209.250 40.500 210.000 ;
        RECT 11.250 208.500 40.500 209.250 ;
        RECT 11.250 207.750 39.750 208.500 ;
        RECT 10.500 207.000 39.750 207.750 ;
        RECT 10.500 205.500 39.000 207.000 ;
        RECT 9.750 204.000 38.250 205.500 ;
        RECT 9.750 203.250 37.500 204.000 ;
        RECT 9.000 202.500 37.500 203.250 ;
        RECT 9.000 201.750 36.750 202.500 ;
        RECT 8.250 201.000 36.750 201.750 ;
        RECT 8.250 199.500 36.000 201.000 ;
        RECT 7.500 197.250 35.250 199.500 ;
        RECT 6.750 195.000 34.500 197.250 ;
        RECT 6.750 194.250 33.750 195.000 ;
        RECT 6.000 193.500 33.750 194.250 ;
        RECT 6.000 192.000 33.000 193.500 ;
        RECT 5.250 191.250 33.000 192.000 ;
        RECT 5.250 189.000 32.250 191.250 ;
        RECT 4.500 186.000 31.500 189.000 ;
        RECT 3.750 183.750 30.750 186.000 ;
        RECT 3.750 182.250 30.000 183.750 ;
        RECT 3.000 180.750 30.000 182.250 ;
        RECT 3.000 178.500 29.250 180.750 ;
        RECT 2.250 177.000 29.250 178.500 ;
        RECT 2.250 174.000 28.500 177.000 ;
        RECT 1.500 173.250 28.500 174.000 ;
        RECT 1.500 168.750 27.750 173.250 ;
        RECT 0.750 168.000 27.750 168.750 ;
        RECT 0.750 161.250 27.000 168.000 ;
        RECT 0.750 159.750 26.250 161.250 ;
        RECT 0.000 143.250 26.250 159.750 ;
        RECT 0.750 141.750 26.250 143.250 ;
        RECT 0.750 134.250 27.000 141.750 ;
        RECT 1.500 129.750 27.750 134.250 ;
        RECT 1.500 129.000 28.500 129.750 ;
        RECT 2.250 126.000 28.500 129.000 ;
        RECT 2.250 124.500 29.250 126.000 ;
        RECT 3.000 122.250 29.250 124.500 ;
        RECT 3.000 120.000 30.000 122.250 ;
        RECT 3.750 119.250 30.000 120.000 ;
        RECT 3.750 117.000 30.750 119.250 ;
        RECT 4.500 114.000 31.500 117.000 ;
        RECT 5.250 111.750 32.250 114.000 ;
        RECT 5.250 111.000 33.000 111.750 ;
        RECT 6.000 109.500 33.000 111.000 ;
        RECT 6.000 108.750 33.750 109.500 ;
        RECT 6.750 108.000 33.750 108.750 ;
        RECT 6.750 105.750 34.500 108.000 ;
        RECT 7.500 103.500 35.250 105.750 ;
        RECT 8.250 102.000 36.000 103.500 ;
        RECT 8.250 101.250 36.750 102.000 ;
        RECT 9.000 100.500 36.750 101.250 ;
        RECT 9.000 99.750 37.500 100.500 ;
        RECT 9.750 99.000 37.500 99.750 ;
        RECT 9.750 97.500 38.250 99.000 ;
        RECT 10.500 96.750 38.250 97.500 ;
        RECT 10.500 95.250 39.000 96.750 ;
        RECT 11.250 93.750 39.750 95.250 ;
        RECT 12.000 92.250 40.500 93.750 ;
        RECT 12.000 91.500 41.250 92.250 ;
        RECT 12.750 90.000 42.000 91.500 ;
        RECT 13.500 88.500 42.750 90.000 ;
        RECT 14.250 87.000 43.500 88.500 ;
        RECT 15.000 86.250 44.250 87.000 ;
        RECT 15.000 85.500 45.000 86.250 ;
        RECT 15.750 84.750 45.000 85.500 ;
        RECT 15.750 84.000 45.750 84.750 ;
        RECT 16.500 82.500 46.500 84.000 ;
        RECT 17.250 81.000 47.250 82.500 ;
        RECT 18.000 80.250 48.000 81.000 ;
        RECT 18.000 79.500 48.750 80.250 ;
        RECT 18.750 78.000 49.500 79.500 ;
        RECT 19.500 77.250 50.250 78.000 ;
        RECT 19.500 76.500 51.000 77.250 ;
        RECT 20.250 75.750 51.000 76.500 ;
        RECT 21.000 75.000 51.750 75.750 ;
        RECT 21.000 74.250 52.500 75.000 ;
        RECT 21.750 73.500 53.250 74.250 ;
        RECT 21.750 72.750 54.000 73.500 ;
        RECT 22.500 72.000 54.000 72.750 ;
        RECT 23.250 71.250 54.750 72.000 ;
        RECT 23.250 70.500 55.500 71.250 ;
        RECT 24.000 69.750 56.250 70.500 ;
        RECT 24.000 69.000 57.000 69.750 ;
        RECT 24.750 68.250 57.750 69.000 ;
        RECT 25.500 67.500 57.750 68.250 ;
        RECT 25.500 66.750 58.500 67.500 ;
        RECT 26.250 66.000 59.250 66.750 ;
        RECT 27.000 65.250 60.000 66.000 ;
        RECT 27.000 64.500 60.750 65.250 ;
        RECT 27.750 63.750 61.500 64.500 ;
        RECT 28.500 63.000 62.250 63.750 ;
        RECT 29.250 62.250 63.000 63.000 ;
        RECT 29.250 61.500 63.750 62.250 ;
        RECT 30.000 60.750 64.500 61.500 ;
        RECT 30.750 60.000 65.250 60.750 ;
        RECT 31.500 59.250 66.000 60.000 ;
        RECT 31.500 58.500 66.750 59.250 ;
        RECT 32.250 57.750 67.500 58.500 ;
        RECT 33.000 57.000 69.000 57.750 ;
        RECT 33.750 56.250 69.750 57.000 ;
        RECT 33.750 55.500 70.500 56.250 ;
        RECT 34.500 54.750 71.250 55.500 ;
        RECT 35.250 54.000 72.000 54.750 ;
        RECT 36.000 53.250 72.750 54.000 ;
        RECT 36.750 52.500 74.250 53.250 ;
        RECT 37.500 51.750 75.000 52.500 ;
        RECT 38.250 51.000 75.750 51.750 ;
        RECT 38.250 50.250 76.500 51.000 ;
        RECT 39.000 49.500 78.000 50.250 ;
        RECT 39.750 48.750 78.750 49.500 ;
        RECT 40.500 48.000 79.500 48.750 ;
        RECT 41.250 47.250 81.000 48.000 ;
        RECT 42.000 46.500 81.750 47.250 ;
        RECT 42.750 45.750 83.250 46.500 ;
        RECT 43.500 45.000 84.000 45.750 ;
        RECT 44.250 44.250 85.500 45.000 ;
        RECT 45.000 43.500 86.250 44.250 ;
        RECT 45.750 42.750 87.750 43.500 ;
        RECT 46.500 42.000 89.250 42.750 ;
        RECT 47.250 41.250 90.750 42.000 ;
        RECT 48.000 40.500 92.250 41.250 ;
        RECT 48.750 39.750 92.250 40.500 ;
        RECT 49.500 39.000 92.250 39.750 ;
        RECT 50.250 38.250 92.250 39.000 ;
        RECT 51.000 37.500 92.250 38.250 ;
        RECT 52.500 36.750 92.250 37.500 ;
        RECT 53.250 36.000 92.250 36.750 ;
        RECT 54.000 35.250 92.250 36.000 ;
        RECT 54.750 34.500 92.250 35.250 ;
        RECT 55.500 33.750 91.500 34.500 ;
        RECT 57.000 33.000 91.500 33.750 ;
        RECT 57.750 32.250 91.500 33.000 ;
        RECT 58.500 31.500 91.500 32.250 ;
        RECT 59.250 30.750 91.500 31.500 ;
        RECT 60.750 30.000 91.500 30.750 ;
        RECT 61.500 29.250 91.500 30.000 ;
        RECT 62.250 28.500 91.500 29.250 ;
        RECT 63.750 27.750 91.500 28.500 ;
        RECT 64.500 27.000 90.750 27.750 ;
        RECT 66.000 26.250 90.750 27.000 ;
        RECT 66.750 25.500 90.750 26.250 ;
        RECT 67.500 24.750 90.750 25.500 ;
        RECT 69.000 24.000 90.750 24.750 ;
        RECT 70.500 23.250 90.750 24.000 ;
        RECT 71.250 22.500 90.750 23.250 ;
        RECT 72.750 21.750 90.750 22.500 ;
        RECT 73.500 21.000 90.000 21.750 ;
        RECT 75.000 20.250 90.000 21.000 ;
        RECT 76.500 19.500 90.000 20.250 ;
        RECT 77.250 18.750 90.000 19.500 ;
        RECT 78.750 18.000 90.000 18.750 ;
        RECT 80.250 17.250 90.000 18.000 ;
        RECT 81.750 16.500 90.000 17.250 ;
        RECT 83.250 15.750 90.000 16.500 ;
        RECT 84.000 15.000 89.250 15.750 ;
        RECT 85.500 14.250 89.250 15.000 ;
        RECT 87.000 13.500 89.250 14.250 ;
        RECT 88.500 12.750 89.250 13.500 ;
    END
  END vss
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER Metal4 ;
        RECT 294.000 438.750 295.500 439.500 ;
        RECT 293.250 438.000 295.500 438.750 ;
        RECT 292.500 436.500 295.500 438.000 ;
        RECT 291.750 435.750 296.250 436.500 ;
        RECT 291.000 435.000 296.250 435.750 ;
        RECT 290.250 434.250 296.250 435.000 ;
        RECT 289.500 433.500 296.250 434.250 ;
        RECT 288.750 432.000 297.000 433.500 ;
        RECT 288.000 431.250 297.000 432.000 ;
        RECT 287.250 430.500 297.750 431.250 ;
        RECT 286.500 429.750 297.750 430.500 ;
        RECT 285.750 428.250 297.750 429.750 ;
        RECT 285.000 427.500 298.500 428.250 ;
        RECT 284.250 426.750 298.500 427.500 ;
        RECT 283.500 426.000 298.500 426.750 ;
        RECT 282.750 425.250 298.500 426.000 ;
        RECT 282.000 423.750 299.250 425.250 ;
        RECT 281.250 423.000 299.250 423.750 ;
        RECT 280.500 422.250 299.250 423.000 ;
        RECT 279.750 421.500 300.000 422.250 ;
        RECT 279.000 420.000 300.000 421.500 ;
        RECT 278.250 419.250 300.000 420.000 ;
        RECT 277.500 418.500 300.750 419.250 ;
        RECT 276.750 417.750 300.750 418.500 ;
        RECT 276.000 416.250 300.750 417.750 ;
        RECT 275.250 415.500 301.500 416.250 ;
        RECT 274.500 414.750 301.500 415.500 ;
        RECT 273.750 414.000 301.500 414.750 ;
        RECT 273.000 413.250 301.500 414.000 ;
        RECT 273.000 412.500 302.250 413.250 ;
        RECT 272.250 411.750 302.250 412.500 ;
        RECT 271.500 411.000 302.250 411.750 ;
        RECT 270.750 410.250 302.250 411.000 ;
        RECT 270.000 409.500 302.250 410.250 ;
        RECT 270.000 408.750 303.000 409.500 ;
        RECT 269.250 408.000 303.000 408.750 ;
        RECT 268.500 407.250 303.000 408.000 ;
        RECT 267.750 406.500 303.000 407.250 ;
        RECT 267.000 405.750 303.000 406.500 ;
        RECT 267.000 405.000 303.750 405.750 ;
        RECT 266.250 404.250 303.750 405.000 ;
        RECT 265.500 403.500 303.750 404.250 ;
        RECT 264.750 402.750 303.750 403.500 ;
        RECT 264.000 402.000 303.750 402.750 ;
        RECT 264.000 401.250 304.500 402.000 ;
        RECT 263.250 400.500 304.500 401.250 ;
        RECT 262.500 399.750 304.500 400.500 ;
        RECT 261.750 399.000 304.500 399.750 ;
        RECT 261.000 397.500 304.500 399.000 ;
        RECT 260.250 396.750 304.500 397.500 ;
        RECT 259.500 396.000 305.250 396.750 ;
        RECT 258.750 395.250 305.250 396.000 ;
        RECT 258.000 393.750 305.250 395.250 ;
        RECT 257.250 393.000 305.250 393.750 ;
        RECT 256.500 392.250 305.250 393.000 ;
        RECT 255.750 390.750 305.250 392.250 ;
        RECT 255.000 390.000 305.250 390.750 ;
        RECT 254.250 389.250 305.250 390.000 ;
        RECT 253.500 388.500 305.250 389.250 ;
        RECT 252.750 387.000 305.250 388.500 ;
        RECT 252.000 386.250 306.000 387.000 ;
        RECT 251.250 385.500 306.000 386.250 ;
        RECT 250.500 384.000 306.000 385.500 ;
        RECT 249.750 383.250 306.000 384.000 ;
        RECT 249.000 382.500 305.250 383.250 ;
        RECT 248.250 381.000 305.250 382.500 ;
        RECT 247.500 380.250 305.250 381.000 ;
        RECT 246.750 379.500 305.250 380.250 ;
        RECT 246.000 378.750 305.250 379.500 ;
        RECT 245.250 377.250 305.250 378.750 ;
        RECT 244.500 376.500 305.250 377.250 ;
        RECT 243.750 375.750 305.250 376.500 ;
        RECT 243.000 374.250 305.250 375.750 ;
        RECT 242.250 373.500 304.500 374.250 ;
        RECT 241.500 372.750 304.500 373.500 ;
        RECT 240.750 371.250 304.500 372.750 ;
        RECT 240.000 370.500 304.500 371.250 ;
        RECT 239.250 369.750 304.500 370.500 ;
        RECT 238.500 368.250 303.750 369.750 ;
        RECT 237.750 367.500 303.750 368.250 ;
        RECT 237.000 366.750 303.750 367.500 ;
        RECT 236.250 365.250 303.750 366.750 ;
        RECT 235.500 364.500 303.000 365.250 ;
        RECT 234.750 363.750 303.000 364.500 ;
        RECT 234.000 362.250 303.000 363.750 ;
        RECT 233.250 361.500 302.250 362.250 ;
        RECT 232.500 360.000 302.250 361.500 ;
        RECT 231.750 359.250 302.250 360.000 ;
        RECT 231.000 358.500 301.500 359.250 ;
        RECT 230.250 357.000 301.500 358.500 ;
        RECT 229.500 356.250 301.500 357.000 ;
        RECT 228.750 355.500 300.750 356.250 ;
        RECT 228.000 354.000 300.750 355.500 ;
        RECT 227.250 353.250 300.750 354.000 ;
        RECT 226.500 351.750 300.000 353.250 ;
        RECT 225.750 351.000 300.000 351.750 ;
        RECT 225.000 350.250 299.250 351.000 ;
        RECT 224.250 348.750 299.250 350.250 ;
        RECT 223.500 348.000 298.500 348.750 ;
        RECT 222.750 346.500 298.500 348.000 ;
        RECT 222.000 345.750 298.500 346.500 ;
        RECT 221.250 345.000 297.750 345.750 ;
        RECT 220.500 343.500 297.750 345.000 ;
        RECT 219.750 342.750 297.000 343.500 ;
        RECT 219.000 341.250 297.000 342.750 ;
        RECT 218.250 340.500 296.250 341.250 ;
        RECT 217.500 339.000 296.250 340.500 ;
        RECT 216.750 338.250 295.500 339.000 ;
        RECT 216.000 336.750 295.500 338.250 ;
        RECT 215.250 336.000 294.750 336.750 ;
        RECT 214.500 335.250 294.750 336.000 ;
        RECT 213.750 334.500 294.750 335.250 ;
        RECT 213.750 333.750 294.000 334.500 ;
        RECT 213.000 333.000 294.000 333.750 ;
        RECT 212.250 332.250 294.000 333.000 ;
        RECT 212.250 331.500 293.250 332.250 ;
        RECT 211.500 330.750 293.250 331.500 ;
        RECT 210.750 330.000 293.250 330.750 ;
        RECT 210.750 329.250 292.500 330.000 ;
        RECT 210.000 328.500 292.500 329.250 ;
        RECT 209.250 327.750 292.500 328.500 ;
        RECT 209.250 327.000 291.750 327.750 ;
        RECT 208.500 326.250 291.750 327.000 ;
        RECT 207.750 325.500 291.750 326.250 ;
        RECT 207.750 324.750 291.000 325.500 ;
        RECT 207.000 324.000 291.000 324.750 ;
        RECT 206.250 322.500 290.250 324.000 ;
        RECT 205.500 321.750 290.250 322.500 ;
        RECT 204.750 320.250 289.500 321.750 ;
        RECT 204.000 319.500 289.500 320.250 ;
        RECT 204.000 318.750 288.750 319.500 ;
        RECT 203.250 318.000 288.750 318.750 ;
        RECT 202.500 316.500 288.000 318.000 ;
        RECT 201.750 315.750 288.000 316.500 ;
        RECT 201.000 314.250 287.250 315.750 ;
        RECT 200.250 313.500 287.250 314.250 ;
        RECT 199.500 312.000 286.500 313.500 ;
        RECT 198.750 310.500 285.750 312.000 ;
        RECT 198.000 309.750 285.750 310.500 ;
        RECT 197.250 308.250 285.000 309.750 ;
        RECT 196.500 307.500 285.000 308.250 ;
        RECT 195.750 306.000 284.250 307.500 ;
        RECT 195.000 304.500 283.500 306.000 ;
        RECT 194.250 303.750 283.500 304.500 ;
        RECT 193.500 302.250 282.750 303.750 ;
        RECT 192.750 300.750 282.000 302.250 ;
        RECT 192.000 300.000 282.000 300.750 ;
        RECT 191.250 298.500 281.250 300.000 ;
        RECT 190.500 297.000 280.500 298.500 ;
        RECT 189.750 296.250 280.500 297.000 ;
        RECT 189.000 294.750 279.750 296.250 ;
        RECT 188.250 293.250 279.000 294.750 ;
        RECT 187.500 292.500 279.000 293.250 ;
        RECT 186.750 291.000 278.250 292.500 ;
        RECT 186.000 289.500 277.500 291.000 ;
        RECT 185.250 288.750 277.500 289.500 ;
        RECT 185.250 288.000 276.750 288.750 ;
        RECT 184.500 287.250 276.750 288.000 ;
        RECT 184.500 286.500 276.000 287.250 ;
        RECT 183.750 285.750 276.000 286.500 ;
        RECT 183.000 285.000 276.000 285.750 ;
        RECT 183.000 284.250 275.250 285.000 ;
        RECT 182.250 283.500 275.250 284.250 ;
        RECT 182.250 282.750 274.500 283.500 ;
        RECT 181.500 282.000 274.500 282.750 ;
        RECT 181.500 281.250 273.750 282.000 ;
        RECT 180.750 279.750 273.750 281.250 ;
        RECT 180.000 279.000 273.000 279.750 ;
        RECT 179.250 278.250 273.000 279.000 ;
        RECT 179.250 277.500 272.250 278.250 ;
        RECT 178.500 276.000 272.250 277.500 ;
        RECT 177.750 274.500 271.500 276.000 ;
        RECT 177.000 273.000 270.750 274.500 ;
        RECT 176.250 271.500 270.000 273.000 ;
        RECT 175.500 270.750 270.000 271.500 ;
        RECT 175.500 270.000 269.250 270.750 ;
        RECT 174.750 269.250 269.250 270.000 ;
        RECT 174.750 268.500 268.500 269.250 ;
        RECT 174.000 267.000 268.500 268.500 ;
        RECT 173.250 265.500 267.750 267.000 ;
        RECT 172.500 264.000 267.000 265.500 ;
        RECT 171.750 262.500 266.250 264.000 ;
        RECT 171.000 261.750 266.250 262.500 ;
        RECT 171.000 261.000 265.500 261.750 ;
        RECT 170.250 260.250 265.500 261.000 ;
        RECT 170.250 259.500 264.750 260.250 ;
        RECT 169.500 258.750 264.750 259.500 ;
        RECT 169.500 258.000 264.000 258.750 ;
        RECT 168.750 256.500 264.000 258.000 ;
        RECT 168.000 255.000 263.250 256.500 ;
        RECT 167.250 253.500 262.500 255.000 ;
        RECT 166.500 252.000 261.750 253.500 ;
        RECT 165.750 251.250 261.750 252.000 ;
        RECT 165.750 250.500 261.000 251.250 ;
        RECT 165.000 249.750 261.000 250.500 ;
        RECT 165.000 248.250 260.250 249.750 ;
        RECT 164.250 246.750 259.500 248.250 ;
        RECT 163.500 246.000 259.500 246.750 ;
        RECT 163.500 245.250 258.750 246.000 ;
        RECT 162.750 244.500 258.750 245.250 ;
        RECT 162.750 243.750 258.000 244.500 ;
        RECT 162.000 243.000 258.000 243.750 ;
        RECT 162.000 241.500 257.250 243.000 ;
        RECT 161.250 240.750 256.500 241.500 ;
        RECT 161.250 240.000 255.750 240.750 ;
        RECT 160.500 239.250 255.000 240.000 ;
        RECT 160.500 238.500 254.250 239.250 ;
        RECT 159.750 237.750 253.500 238.500 ;
        RECT 159.750 237.000 252.750 237.750 ;
        RECT 159.000 236.250 252.000 237.000 ;
        RECT 159.000 235.500 251.250 236.250 ;
        RECT 159.000 234.750 250.500 235.500 ;
        RECT 158.250 234.000 249.750 234.750 ;
        RECT 158.250 233.250 249.000 234.000 ;
        RECT 157.500 232.500 248.250 233.250 ;
        RECT 157.500 231.750 247.500 232.500 ;
        RECT 157.500 231.000 246.750 231.750 ;
        RECT 156.750 230.250 246.000 231.000 ;
        RECT 156.750 229.500 245.250 230.250 ;
        RECT 156.000 228.750 244.500 229.500 ;
        RECT 156.000 228.000 243.750 228.750 ;
        RECT 155.250 227.250 243.000 228.000 ;
        RECT 155.250 226.500 242.250 227.250 ;
        RECT 155.250 225.750 241.500 226.500 ;
        RECT 154.500 224.250 240.750 225.750 ;
        RECT 153.750 223.500 240.000 224.250 ;
        RECT 153.750 222.750 239.250 223.500 ;
        RECT 153.750 222.000 238.500 222.750 ;
        RECT 153.000 221.250 237.750 222.000 ;
        RECT 153.000 220.500 237.000 221.250 ;
        RECT 152.250 219.750 236.250 220.500 ;
        RECT 152.250 219.000 235.500 219.750 ;
        RECT 152.250 218.250 234.750 219.000 ;
        RECT 151.500 217.500 234.000 218.250 ;
        RECT 151.500 216.750 233.250 217.500 ;
        RECT 150.750 216.000 232.500 216.750 ;
        RECT 150.750 215.250 231.750 216.000 ;
        RECT 150.750 214.500 231.000 215.250 ;
        RECT 150.000 213.750 230.250 214.500 ;
        RECT 150.000 213.000 229.500 213.750 ;
        RECT 149.250 212.250 228.750 213.000 ;
        RECT 149.250 211.500 228.000 212.250 ;
        RECT 149.250 210.750 227.250 211.500 ;
        RECT 148.500 210.000 226.500 210.750 ;
        RECT 148.500 209.250 225.750 210.000 ;
        RECT 148.500 208.500 225.000 209.250 ;
        RECT 147.750 207.750 224.250 208.500 ;
        RECT 147.750 207.000 223.500 207.750 ;
        RECT 147.000 206.250 222.750 207.000 ;
        RECT 147.000 205.500 222.000 206.250 ;
        RECT 147.000 204.750 221.250 205.500 ;
        RECT 146.250 204.000 220.500 204.750 ;
        RECT 146.250 203.250 219.750 204.000 ;
        RECT 146.250 202.500 219.000 203.250 ;
        RECT 145.500 201.750 219.000 202.500 ;
        RECT 145.500 201.000 218.250 201.750 ;
        RECT 144.750 200.250 217.500 201.000 ;
        RECT 144.750 199.500 216.750 200.250 ;
        RECT 144.750 198.750 216.000 199.500 ;
        RECT 144.000 198.000 215.250 198.750 ;
        RECT 144.000 197.250 214.500 198.000 ;
        RECT 144.000 196.500 213.750 197.250 ;
        RECT 143.250 195.750 213.000 196.500 ;
        RECT 143.250 195.000 212.250 195.750 ;
        RECT 143.250 194.250 211.500 195.000 ;
        RECT 142.500 193.500 210.750 194.250 ;
        RECT 142.500 192.750 210.000 193.500 ;
        RECT 141.750 191.250 209.250 192.750 ;
        RECT 141.750 190.500 208.500 191.250 ;
        RECT 141.000 189.750 207.750 190.500 ;
        RECT 141.000 189.000 207.000 189.750 ;
        RECT 141.000 188.250 206.250 189.000 ;
        RECT 140.250 187.500 205.500 188.250 ;
        RECT 140.250 186.750 204.750 187.500 ;
        RECT 140.250 186.000 204.000 186.750 ;
        RECT 139.500 185.250 204.000 186.000 ;
        RECT 139.500 184.500 203.250 185.250 ;
        RECT 139.500 183.750 202.500 184.500 ;
        RECT 138.750 183.000 201.750 183.750 ;
        RECT 138.750 182.250 201.000 183.000 ;
        RECT 138.750 181.500 200.250 182.250 ;
        RECT 138.000 180.000 199.500 181.500 ;
        RECT 138.000 179.250 198.750 180.000 ;
        RECT 137.250 178.500 198.000 179.250 ;
        RECT 137.250 177.750 197.250 178.500 ;
        RECT 137.250 177.000 196.500 177.750 ;
        RECT 136.500 175.500 195.750 177.000 ;
        RECT 136.500 174.750 195.000 175.500 ;
        RECT 135.750 174.000 194.250 174.750 ;
        RECT 135.750 173.250 193.500 174.000 ;
        RECT 135.750 172.500 192.750 173.250 ;
        RECT 135.000 171.000 192.000 172.500 ;
        RECT 135.000 170.250 191.250 171.000 ;
        RECT 134.250 169.500 190.500 170.250 ;
        RECT 134.250 168.750 189.750 169.500 ;
        RECT 134.250 167.250 189.000 168.750 ;
        RECT 133.500 166.500 188.250 167.250 ;
        RECT 133.500 165.750 187.500 166.500 ;
        RECT 133.500 165.000 186.750 165.750 ;
        RECT 132.750 164.250 186.750 165.000 ;
        RECT 132.750 163.500 186.000 164.250 ;
        RECT 132.750 162.750 185.250 163.500 ;
        RECT 132.000 162.000 184.500 162.750 ;
        RECT 132.000 160.500 183.750 162.000 ;
        RECT 131.250 159.750 183.000 160.500 ;
        RECT 131.250 159.000 182.250 159.750 ;
        RECT 131.250 158.250 181.500 159.000 ;
        RECT 130.500 157.500 181.500 158.250 ;
        RECT 130.500 156.750 180.750 157.500 ;
        RECT 130.500 156.000 180.000 156.750 ;
        RECT 130.500 155.250 179.250 156.000 ;
        RECT 129.750 154.500 179.250 155.250 ;
        RECT 129.750 153.750 178.500 154.500 ;
        RECT 129.750 153.000 177.750 153.750 ;
        RECT 129.000 151.500 177.000 153.000 ;
        RECT 129.000 150.750 176.250 151.500 ;
        RECT 128.250 150.000 175.500 150.750 ;
        RECT 128.250 148.500 174.750 150.000 ;
        RECT 128.250 147.750 174.000 148.500 ;
        RECT 127.500 146.250 173.250 147.750 ;
        RECT 127.500 145.500 172.500 146.250 ;
        RECT 126.750 144.750 171.750 145.500 ;
        RECT 126.750 143.250 171.000 144.750 ;
        RECT 126.750 142.500 170.250 143.250 ;
        RECT 126.000 141.750 169.500 142.500 ;
        RECT 126.000 140.250 168.750 141.750 ;
        RECT 125.250 139.500 168.000 140.250 ;
        RECT 125.250 138.000 167.250 139.500 ;
        RECT 124.500 137.250 166.500 138.000 ;
        RECT 124.500 136.500 165.750 137.250 ;
        RECT 124.500 135.000 165.000 136.500 ;
        RECT 123.750 134.250 164.250 135.000 ;
        RECT 123.750 133.500 163.500 134.250 ;
        RECT 123.750 132.750 162.750 133.500 ;
        RECT 123.000 132.000 162.750 132.750 ;
        RECT 123.000 131.250 162.000 132.000 ;
        RECT 123.000 129.750 161.250 131.250 ;
        RECT 122.250 129.000 160.500 129.750 ;
        RECT 122.250 127.500 159.750 129.000 ;
        RECT 121.500 126.750 159.000 127.500 ;
        RECT 121.500 126.000 158.250 126.750 ;
        RECT 121.500 124.500 157.500 126.000 ;
        RECT 120.750 123.750 156.750 124.500 ;
        RECT 120.750 122.250 156.000 123.750 ;
        RECT 120.000 121.500 155.250 122.250 ;
        RECT 120.000 120.000 154.500 121.500 ;
        RECT 120.000 119.250 153.750 120.000 ;
        RECT 119.250 117.750 153.000 119.250 ;
        RECT 119.250 117.000 152.250 117.750 ;
        RECT 118.500 115.500 151.500 117.000 ;
        RECT 118.500 114.750 150.750 115.500 ;
        RECT 118.500 114.000 150.000 114.750 ;
        RECT 117.750 113.250 150.000 114.000 ;
        RECT 117.750 112.500 149.250 113.250 ;
        RECT 117.750 111.750 148.500 112.500 ;
        RECT 117.000 111.000 148.500 111.750 ;
        RECT 117.000 110.250 147.750 111.000 ;
        RECT 117.000 108.750 147.000 110.250 ;
        RECT 116.250 108.000 146.250 108.750 ;
        RECT 116.250 106.500 145.500 108.000 ;
        RECT 115.500 105.750 144.750 106.500 ;
        RECT 115.500 104.250 144.000 105.750 ;
        RECT 115.500 103.500 143.250 104.250 ;
        RECT 114.750 102.000 142.500 103.500 ;
        RECT 114.750 101.250 141.750 102.000 ;
        RECT 114.750 100.500 141.000 101.250 ;
        RECT 114.000 99.750 141.000 100.500 ;
        RECT 114.000 98.250 140.250 99.750 ;
        RECT 114.000 97.500 139.500 98.250 ;
        RECT 113.250 96.000 138.750 97.500 ;
        RECT 113.250 95.250 138.000 96.000 ;
        RECT 112.500 94.500 138.000 95.250 ;
        RECT 112.500 93.750 137.250 94.500 ;
        RECT 112.500 92.250 136.500 93.750 ;
        RECT 111.750 91.500 135.750 92.250 ;
        RECT 111.750 90.000 135.000 91.500 ;
        RECT 111.750 89.250 134.250 90.000 ;
        RECT 111.000 88.500 134.250 89.250 ;
        RECT 111.000 87.000 133.500 88.500 ;
        RECT 111.000 86.250 132.750 87.000 ;
        RECT 110.250 84.750 132.000 86.250 ;
        RECT 110.250 83.250 131.250 84.750 ;
        RECT 109.500 81.750 130.500 83.250 ;
        RECT 109.500 81.000 129.750 81.750 ;
        RECT 109.500 80.250 129.000 81.000 ;
        RECT 108.750 79.500 129.000 80.250 ;
        RECT 108.750 78.000 128.250 79.500 ;
        RECT 108.750 77.250 127.500 78.000 ;
        RECT 108.000 76.500 127.500 77.250 ;
        RECT 108.000 75.000 126.750 76.500 ;
        RECT 108.000 73.500 126.000 75.000 ;
        RECT 107.250 72.750 125.250 73.500 ;
        RECT 107.250 71.250 124.500 72.750 ;
        RECT 107.250 70.500 123.750 71.250 ;
        RECT 106.500 69.750 123.750 70.500 ;
        RECT 106.500 68.250 123.000 69.750 ;
        RECT 106.500 66.750 122.250 68.250 ;
        RECT 105.750 65.250 121.500 66.750 ;
        RECT 105.750 63.750 120.750 65.250 ;
        RECT 105.000 62.250 120.000 63.750 ;
        RECT 105.000 60.750 119.250 62.250 ;
        RECT 105.000 60.000 118.500 60.750 ;
        RECT 104.250 59.250 118.500 60.000 ;
        RECT 104.250 57.750 117.750 59.250 ;
        RECT 104.250 56.250 117.000 57.750 ;
        RECT 103.500 54.750 116.250 56.250 ;
        RECT 103.500 53.250 115.500 54.750 ;
        RECT 103.500 52.500 114.750 53.250 ;
        RECT 102.750 51.750 114.750 52.500 ;
        RECT 102.750 50.250 114.000 51.750 ;
        RECT 102.750 49.500 113.250 50.250 ;
        RECT 102.000 48.750 113.250 49.500 ;
        RECT 102.000 47.250 112.500 48.750 ;
        RECT 102.000 45.750 111.750 47.250 ;
        RECT 101.250 44.250 111.000 45.750 ;
        RECT 101.250 42.750 110.250 44.250 ;
        RECT 101.250 41.250 109.500 42.750 ;
        RECT 100.500 39.750 108.750 41.250 ;
        RECT 100.500 38.250 108.000 39.750 ;
        RECT 100.500 37.500 107.250 38.250 ;
        RECT 99.750 36.750 107.250 37.500 ;
        RECT 99.750 35.250 106.500 36.750 ;
        RECT 99.750 33.750 105.750 35.250 ;
        RECT 99.000 32.250 105.000 33.750 ;
        RECT 99.000 30.750 104.250 32.250 ;
        RECT 99.000 30.000 103.500 30.750 ;
        RECT 98.250 29.250 103.500 30.000 ;
        RECT 98.250 27.750 102.750 29.250 ;
        RECT 98.250 26.250 102.000 27.750 ;
        RECT 97.500 25.500 102.000 26.250 ;
        RECT 97.500 24.000 101.250 25.500 ;
        RECT 97.500 22.500 100.500 24.000 ;
        RECT 97.500 21.750 99.750 22.500 ;
        RECT 96.750 21.000 99.750 21.750 ;
        RECT 96.750 19.500 99.000 21.000 ;
        RECT 96.750 18.000 98.250 19.500 ;
        RECT 96.000 16.500 97.500 18.000 ;
        RECT 96.000 15.000 96.750 16.500 ;
    END
  END vdd
  OBS
      LAYER Metal2 ;
        RECT 0.000 0.000 375.000 440.250 ;
      LAYER Metal3 ;
        RECT 0.000 0.000 375.000 440.250 ;
      LAYER Metal4 ;
        RECT 365.250 313.500 366.000 314.250 ;
        RECT 364.500 312.750 366.000 313.500 ;
        RECT 363.000 312.000 366.000 312.750 ;
        RECT 362.250 311.250 366.000 312.000 ;
        RECT 360.750 310.500 366.000 311.250 ;
        RECT 360.000 309.750 366.000 310.500 ;
        RECT 358.500 309.000 366.000 309.750 ;
        RECT 357.750 308.250 366.000 309.000 ;
        RECT 356.250 307.500 366.000 308.250 ;
        RECT 354.750 306.750 366.000 307.500 ;
        RECT 354.000 306.000 366.000 306.750 ;
        RECT 352.500 305.250 366.000 306.000 ;
        RECT 351.750 304.500 366.000 305.250 ;
        RECT 350.250 303.750 366.000 304.500 ;
        RECT 349.500 303.000 366.000 303.750 ;
        RECT 348.000 302.250 366.000 303.000 ;
        RECT 347.250 301.500 366.000 302.250 ;
        RECT 345.750 300.750 366.000 301.500 ;
        RECT 345.000 300.000 366.000 300.750 ;
        RECT 343.500 299.250 366.000 300.000 ;
        RECT 342.750 298.500 366.000 299.250 ;
        RECT 341.250 297.750 366.000 298.500 ;
        RECT 340.500 297.000 366.000 297.750 ;
        RECT 339.000 296.250 366.000 297.000 ;
        RECT 338.250 295.500 366.000 296.250 ;
        RECT 337.500 294.750 366.000 295.500 ;
        RECT 336.000 294.000 366.000 294.750 ;
        RECT 335.250 293.250 366.000 294.000 ;
        RECT 333.750 292.500 366.000 293.250 ;
        RECT 333.000 291.750 366.000 292.500 ;
        RECT 331.500 291.000 366.000 291.750 ;
        RECT 330.750 290.250 366.000 291.000 ;
        RECT 330.000 289.500 366.000 290.250 ;
        RECT 328.500 288.750 366.000 289.500 ;
        RECT 327.750 288.000 366.000 288.750 ;
        RECT 326.250 287.250 366.000 288.000 ;
        RECT 325.500 286.500 366.000 287.250 ;
        RECT 324.750 285.750 366.000 286.500 ;
        RECT 323.250 285.000 366.000 285.750 ;
        RECT 322.500 284.250 366.000 285.000 ;
        RECT 321.750 283.500 366.000 284.250 ;
        RECT 320.250 282.750 365.250 283.500 ;
        RECT 319.500 282.000 365.250 282.750 ;
        RECT 318.750 281.250 365.250 282.000 ;
        RECT 317.250 280.500 365.250 281.250 ;
        RECT 316.500 279.750 365.250 280.500 ;
        RECT 315.750 279.000 365.250 279.750 ;
        RECT 314.250 278.250 365.250 279.000 ;
        RECT 313.500 277.500 365.250 278.250 ;
        RECT 312.750 276.750 364.500 277.500 ;
        RECT 311.250 276.000 364.500 276.750 ;
        RECT 310.500 275.250 364.500 276.000 ;
        RECT 309.750 274.500 364.500 275.250 ;
        RECT 308.250 273.750 364.500 274.500 ;
        RECT 307.500 273.000 363.750 273.750 ;
        RECT 306.750 272.250 363.750 273.000 ;
        RECT 306.000 271.500 363.750 272.250 ;
        RECT 304.500 270.750 363.750 271.500 ;
        RECT 303.750 270.000 363.000 270.750 ;
        RECT 303.000 269.250 363.000 270.000 ;
        RECT 301.500 268.500 363.000 269.250 ;
        RECT 300.750 267.750 363.000 268.500 ;
        RECT 300.000 267.000 362.250 267.750 ;
        RECT 299.250 266.250 362.250 267.000 ;
        RECT 298.500 265.500 362.250 266.250 ;
        RECT 297.000 264.750 362.250 265.500 ;
        RECT 296.250 264.000 361.500 264.750 ;
        RECT 295.500 263.250 361.500 264.000 ;
        RECT 294.750 262.500 360.750 263.250 ;
        RECT 293.250 261.750 360.750 262.500 ;
        RECT 292.500 261.000 360.000 261.750 ;
        RECT 291.750 260.250 360.000 261.000 ;
        RECT 291.000 259.500 360.000 260.250 ;
        RECT 289.500 258.750 359.250 259.500 ;
        RECT 288.750 258.000 359.250 258.750 ;
        RECT 288.000 257.250 358.500 258.000 ;
        RECT 287.250 256.500 358.500 257.250 ;
        RECT 286.500 255.750 357.750 256.500 ;
        RECT 285.000 255.000 357.750 255.750 ;
        RECT 284.250 254.250 357.750 255.000 ;
        RECT 283.500 253.500 357.000 254.250 ;
        RECT 282.750 252.750 357.000 253.500 ;
        RECT 282.000 252.000 356.250 252.750 ;
        RECT 281.250 251.250 355.500 252.000 ;
        RECT 279.750 250.500 355.500 251.250 ;
        RECT 279.000 249.750 354.750 250.500 ;
        RECT 278.250 249.000 354.750 249.750 ;
        RECT 277.500 248.250 354.000 249.000 ;
        RECT 276.750 247.500 353.250 248.250 ;
        RECT 275.250 246.750 353.250 247.500 ;
        RECT 274.500 246.000 352.500 246.750 ;
        RECT 273.750 245.250 352.500 246.000 ;
        RECT 273.000 244.500 351.750 245.250 ;
        RECT 272.250 243.750 351.000 244.500 ;
        RECT 271.500 243.000 351.000 243.750 ;
        RECT 270.750 242.250 350.250 243.000 ;
        RECT 270.000 241.500 350.250 242.250 ;
        RECT 268.500 240.750 349.500 241.500 ;
        RECT 267.750 240.000 348.750 240.750 ;
        RECT 267.000 239.250 348.750 240.000 ;
        RECT 266.250 238.500 348.000 239.250 ;
        RECT 265.500 237.750 347.250 238.500 ;
        RECT 264.750 237.000 347.250 237.750 ;
        RECT 264.000 236.250 346.500 237.000 ;
        RECT 263.250 235.500 345.750 236.250 ;
        RECT 261.750 234.750 345.000 235.500 ;
        RECT 261.000 234.000 345.000 234.750 ;
        RECT 260.250 233.250 344.250 234.000 ;
        RECT 259.500 232.500 343.500 233.250 ;
        RECT 258.750 231.750 343.500 232.500 ;
        RECT 258.000 231.000 342.750 231.750 ;
        RECT 257.250 230.250 342.000 231.000 ;
        RECT 256.500 229.500 341.250 230.250 ;
        RECT 255.750 228.750 341.250 229.500 ;
        RECT 255.000 228.000 340.500 228.750 ;
        RECT 254.250 227.250 339.750 228.000 ;
        RECT 252.750 226.500 339.750 227.250 ;
        RECT 252.000 225.750 339.000 226.500 ;
        RECT 251.250 225.000 338.250 225.750 ;
        RECT 250.500 224.250 337.500 225.000 ;
        RECT 249.750 223.500 336.750 224.250 ;
        RECT 249.000 222.750 336.750 223.500 ;
        RECT 248.250 222.000 336.000 222.750 ;
        RECT 247.500 221.250 335.250 222.000 ;
        RECT 246.750 220.500 334.500 221.250 ;
        RECT 246.000 219.750 334.500 220.500 ;
        RECT 245.250 219.000 333.750 219.750 ;
        RECT 244.500 218.250 333.000 219.000 ;
        RECT 243.750 217.500 332.250 218.250 ;
        RECT 243.000 216.750 331.500 217.500 ;
        RECT 242.250 216.000 331.500 216.750 ;
        RECT 241.500 215.250 330.750 216.000 ;
        RECT 240.750 214.500 330.000 215.250 ;
        RECT 240.000 213.750 329.250 214.500 ;
        RECT 238.500 213.000 329.250 213.750 ;
        RECT 237.750 212.250 328.500 213.000 ;
        RECT 237.000 211.500 327.750 212.250 ;
        RECT 236.250 210.750 327.000 211.500 ;
        RECT 235.500 210.000 326.250 210.750 ;
        RECT 234.750 209.250 326.250 210.000 ;
        RECT 234.000 208.500 325.500 209.250 ;
        RECT 233.250 207.750 324.750 208.500 ;
        RECT 232.500 207.000 324.000 207.750 ;
        RECT 231.750 206.250 323.250 207.000 ;
        RECT 231.000 205.500 323.250 206.250 ;
        RECT 230.250 204.750 322.500 205.500 ;
        RECT 229.500 204.000 321.750 204.750 ;
        RECT 228.750 203.250 321.000 204.000 ;
        RECT 228.000 202.500 320.250 203.250 ;
        RECT 227.250 201.750 320.250 202.500 ;
        RECT 226.500 201.000 319.500 201.750 ;
        RECT 225.750 200.250 318.750 201.000 ;
        RECT 225.000 199.500 318.000 200.250 ;
        RECT 224.250 198.750 317.250 199.500 ;
        RECT 223.500 198.000 316.500 198.750 ;
        RECT 222.750 197.250 316.500 198.000 ;
        RECT 222.000 196.500 315.750 197.250 ;
        RECT 221.250 195.750 315.000 196.500 ;
        RECT 220.500 195.000 314.250 195.750 ;
        RECT 219.750 194.250 313.500 195.000 ;
        RECT 219.000 193.500 313.500 194.250 ;
        RECT 218.250 192.750 312.750 193.500 ;
        RECT 217.500 192.000 312.000 192.750 ;
        RECT 216.750 191.250 311.250 192.000 ;
        RECT 216.750 190.500 310.500 191.250 ;
        RECT 216.000 189.750 310.500 190.500 ;
        RECT 215.250 189.000 309.750 189.750 ;
        RECT 214.500 188.250 309.000 189.000 ;
        RECT 213.750 187.500 308.250 188.250 ;
        RECT 213.000 186.750 307.500 187.500 ;
        RECT 212.250 186.000 307.500 186.750 ;
        RECT 211.500 185.250 306.750 186.000 ;
        RECT 210.750 184.500 306.000 185.250 ;
        RECT 210.000 183.750 305.250 184.500 ;
        RECT 209.250 183.000 304.500 183.750 ;
        RECT 208.500 182.250 303.750 183.000 ;
        RECT 207.750 181.500 303.750 182.250 ;
        RECT 207.000 180.750 303.000 181.500 ;
        RECT 206.250 180.000 302.250 180.750 ;
        RECT 206.250 179.250 301.500 180.000 ;
        RECT 205.500 178.500 300.750 179.250 ;
        RECT 204.750 177.750 300.750 178.500 ;
        RECT 204.000 177.000 300.000 177.750 ;
        RECT 203.250 176.250 299.250 177.000 ;
        RECT 202.500 175.500 298.500 176.250 ;
        RECT 201.750 174.750 297.750 175.500 ;
        RECT 201.000 174.000 297.750 174.750 ;
        RECT 200.250 173.250 297.000 174.000 ;
        RECT 200.250 172.500 296.250 173.250 ;
        RECT 199.500 171.750 295.500 172.500 ;
        RECT 198.750 171.000 294.750 171.750 ;
        RECT 198.000 170.250 294.000 171.000 ;
        RECT 197.250 169.500 294.000 170.250 ;
        RECT 301.500 169.500 302.250 170.250 ;
        RECT 196.500 168.750 293.250 169.500 ;
        RECT 300.750 168.750 302.250 169.500 ;
        RECT 196.500 168.000 292.500 168.750 ;
        RECT 300.000 168.000 303.000 168.750 ;
        RECT 195.750 167.250 291.750 168.000 ;
        RECT 299.250 167.250 303.000 168.000 ;
        RECT 195.000 166.500 291.000 167.250 ;
        RECT 298.500 166.500 303.000 167.250 ;
        RECT 194.250 165.750 291.000 166.500 ;
        RECT 193.500 165.000 290.250 165.750 ;
        RECT 297.750 165.000 303.000 166.500 ;
        RECT 192.750 164.250 289.500 165.000 ;
        RECT 297.000 164.250 303.000 165.000 ;
        RECT 192.750 163.500 288.750 164.250 ;
        RECT 296.250 163.500 303.750 164.250 ;
        RECT 192.000 162.750 288.000 163.500 ;
        RECT 295.500 162.750 303.750 163.500 ;
        RECT 191.250 162.000 287.250 162.750 ;
        RECT 294.750 162.000 303.750 162.750 ;
        RECT 190.500 161.250 287.250 162.000 ;
        RECT 294.000 161.250 303.750 162.000 ;
        RECT 189.750 160.500 286.500 161.250 ;
        RECT 189.750 159.750 285.750 160.500 ;
        RECT 293.250 159.750 303.750 161.250 ;
        RECT 189.000 159.000 285.000 159.750 ;
        RECT 292.500 159.000 303.750 159.750 ;
        RECT 188.250 158.250 284.250 159.000 ;
        RECT 291.750 158.250 303.750 159.000 ;
        RECT 187.500 157.500 284.250 158.250 ;
        RECT 291.000 157.500 303.750 158.250 ;
        RECT 187.500 156.750 283.500 157.500 ;
        RECT 290.250 156.750 303.750 157.500 ;
        RECT 186.750 156.000 282.750 156.750 ;
        RECT 289.500 156.000 303.750 156.750 ;
        RECT 186.000 155.250 282.000 156.000 ;
        RECT 288.750 155.250 303.750 156.000 ;
        RECT 185.250 154.500 281.250 155.250 ;
        RECT 184.500 153.750 281.250 154.500 ;
        RECT 288.000 153.750 303.750 155.250 ;
        RECT 184.500 153.000 280.500 153.750 ;
        RECT 287.250 153.000 303.750 153.750 ;
        RECT 183.750 152.250 279.750 153.000 ;
        RECT 286.500 152.250 303.750 153.000 ;
        RECT 183.000 151.500 279.000 152.250 ;
        RECT 285.750 151.500 303.750 152.250 ;
        RECT 182.250 150.750 278.250 151.500 ;
        RECT 285.000 150.750 303.750 151.500 ;
        RECT 182.250 150.000 277.500 150.750 ;
        RECT 284.250 150.000 303.750 150.750 ;
        RECT 181.500 149.250 277.500 150.000 ;
        RECT 283.500 149.250 303.750 150.000 ;
        RECT 372.000 149.250 375.000 150.000 ;
        RECT 180.750 148.500 276.750 149.250 ;
        RECT 180.750 147.750 276.000 148.500 ;
        RECT 282.750 147.750 303.750 149.250 ;
        RECT 369.000 148.500 374.250 149.250 ;
        RECT 366.000 147.750 374.250 148.500 ;
        RECT 180.000 147.000 275.250 147.750 ;
        RECT 282.000 147.000 303.750 147.750 ;
        RECT 363.000 147.000 373.500 147.750 ;
        RECT 179.250 146.250 274.500 147.000 ;
        RECT 281.250 146.250 303.750 147.000 ;
        RECT 359.250 146.250 373.500 147.000 ;
        RECT 178.500 145.500 274.500 146.250 ;
        RECT 280.500 145.500 303.750 146.250 ;
        RECT 356.250 145.500 373.500 146.250 ;
        RECT 178.500 144.750 273.750 145.500 ;
        RECT 279.750 144.750 303.750 145.500 ;
        RECT 353.250 144.750 372.750 145.500 ;
        RECT 177.750 144.000 273.000 144.750 ;
        RECT 279.000 144.000 303.750 144.750 ;
        RECT 350.250 144.000 372.750 144.750 ;
        RECT 177.000 143.250 272.250 144.000 ;
        RECT 278.250 143.250 303.750 144.000 ;
        RECT 347.250 143.250 372.000 144.000 ;
        RECT 176.250 142.500 271.500 143.250 ;
        RECT 278.250 142.500 303.000 143.250 ;
        RECT 344.250 142.500 372.000 143.250 ;
        RECT 176.250 141.750 270.750 142.500 ;
        RECT 277.500 141.750 303.000 142.500 ;
        RECT 341.250 141.750 372.000 142.500 ;
        RECT 175.500 141.000 270.750 141.750 ;
        RECT 276.750 141.000 303.000 141.750 ;
        RECT 338.250 141.000 371.250 141.750 ;
        RECT 174.750 140.250 270.000 141.000 ;
        RECT 276.000 140.250 303.000 141.000 ;
        RECT 335.250 140.250 371.250 141.000 ;
        RECT 174.750 139.500 269.250 140.250 ;
        RECT 276.000 139.500 301.500 140.250 ;
        RECT 332.250 139.500 370.500 140.250 ;
        RECT 174.000 138.750 268.500 139.500 ;
        RECT 276.000 138.750 299.250 139.500 ;
        RECT 329.250 138.750 370.500 139.500 ;
        RECT 173.250 137.250 267.750 138.750 ;
        RECT 276.000 138.000 297.750 138.750 ;
        RECT 326.250 138.000 369.750 138.750 ;
        RECT 276.000 137.250 295.500 138.000 ;
        RECT 324.000 137.250 369.750 138.000 ;
        RECT 172.500 136.500 267.000 137.250 ;
        RECT 276.000 136.500 293.250 137.250 ;
        RECT 321.000 136.500 369.000 137.250 ;
        RECT 171.750 135.750 266.250 136.500 ;
        RECT 276.000 135.750 291.750 136.500 ;
        RECT 318.000 135.750 369.000 136.500 ;
        RECT 171.000 135.000 265.500 135.750 ;
        RECT 276.000 135.000 289.500 135.750 ;
        RECT 315.000 135.000 368.250 135.750 ;
        RECT 171.000 134.250 264.750 135.000 ;
        RECT 276.000 134.250 287.250 135.000 ;
        RECT 312.750 134.250 368.250 135.000 ;
        RECT 170.250 133.500 264.000 134.250 ;
        RECT 169.500 132.750 264.000 133.500 ;
        RECT 276.000 133.500 285.000 134.250 ;
        RECT 309.750 133.500 367.500 134.250 ;
        RECT 276.000 132.750 283.500 133.500 ;
        RECT 306.750 132.750 367.500 133.500 ;
        RECT 169.500 132.000 263.250 132.750 ;
        RECT 276.000 132.000 281.250 132.750 ;
        RECT 304.500 132.000 366.750 132.750 ;
        RECT 168.750 131.250 262.500 132.000 ;
        RECT 276.000 131.250 279.000 132.000 ;
        RECT 301.500 131.250 366.750 132.000 ;
        RECT 168.000 130.500 261.750 131.250 ;
        RECT 275.250 130.500 276.750 131.250 ;
        RECT 299.250 130.500 366.000 131.250 ;
        RECT 168.000 129.750 261.000 130.500 ;
        RECT 296.250 129.750 365.250 130.500 ;
        RECT 167.250 129.000 260.250 129.750 ;
        RECT 294.000 129.000 365.250 129.750 ;
        RECT 166.500 128.250 258.750 129.000 ;
        RECT 291.000 128.250 364.500 129.000 ;
        RECT 166.500 127.500 257.250 128.250 ;
        RECT 288.750 127.500 364.500 128.250 ;
        RECT 165.750 126.750 255.750 127.500 ;
        RECT 285.750 126.750 363.750 127.500 ;
        RECT 165.000 126.000 254.250 126.750 ;
        RECT 283.500 126.000 363.000 126.750 ;
        RECT 165.000 125.250 252.750 126.000 ;
        RECT 281.250 125.250 362.250 126.000 ;
        RECT 164.250 124.500 251.250 125.250 ;
        RECT 279.000 124.500 361.500 125.250 ;
        RECT 163.500 123.750 249.750 124.500 ;
        RECT 276.750 123.750 361.500 124.500 ;
        RECT 163.500 123.000 248.250 123.750 ;
        RECT 274.500 123.000 360.750 123.750 ;
        RECT 162.750 122.250 246.750 123.000 ;
        RECT 272.250 122.250 360.000 123.000 ;
        RECT 162.000 121.500 245.250 122.250 ;
        RECT 270.000 121.500 359.250 122.250 ;
        RECT 162.000 120.750 243.750 121.500 ;
        RECT 267.750 120.750 358.500 121.500 ;
        RECT 161.250 120.000 242.250 120.750 ;
        RECT 265.500 120.000 357.750 120.750 ;
        RECT 160.500 119.250 240.750 120.000 ;
        RECT 263.250 119.250 357.750 120.000 ;
        RECT 160.500 118.500 240.000 119.250 ;
        RECT 261.750 118.500 357.000 119.250 ;
        RECT 159.750 117.750 238.500 118.500 ;
        RECT 259.500 117.750 356.250 118.500 ;
        RECT 159.000 117.000 237.000 117.750 ;
        RECT 257.250 117.000 355.500 117.750 ;
        RECT 159.000 116.250 235.500 117.000 ;
        RECT 255.750 116.250 354.750 117.000 ;
        RECT 158.250 115.500 234.000 116.250 ;
        RECT 253.500 115.500 354.000 116.250 ;
        RECT 157.500 114.750 232.500 115.500 ;
        RECT 252.000 114.750 353.250 115.500 ;
        RECT 157.500 114.000 231.000 114.750 ;
        RECT 249.750 114.000 352.500 114.750 ;
        RECT 156.750 113.250 229.500 114.000 ;
        RECT 248.250 113.250 351.000 114.000 ;
        RECT 156.000 112.500 228.750 113.250 ;
        RECT 246.000 112.500 350.250 113.250 ;
        RECT 156.000 111.750 227.250 112.500 ;
        RECT 244.500 111.750 349.500 112.500 ;
        RECT 155.250 111.000 225.750 111.750 ;
        RECT 243.000 111.000 348.750 111.750 ;
        RECT 154.500 110.250 224.250 111.000 ;
        RECT 241.500 110.250 348.000 111.000 ;
        RECT 154.500 109.500 222.750 110.250 ;
        RECT 240.000 109.500 346.500 110.250 ;
        RECT 153.750 108.750 221.250 109.500 ;
        RECT 237.750 108.750 345.750 109.500 ;
        RECT 153.000 108.000 220.500 108.750 ;
        RECT 236.250 108.000 345.000 108.750 ;
        RECT 153.000 107.250 219.000 108.000 ;
        RECT 234.750 107.250 344.250 108.000 ;
        RECT 152.250 106.500 217.500 107.250 ;
        RECT 233.250 106.500 342.750 107.250 ;
        RECT 152.250 105.750 216.000 106.500 ;
        RECT 231.750 105.750 342.000 106.500 ;
        RECT 151.500 105.000 214.500 105.750 ;
        RECT 230.250 105.000 341.250 105.750 ;
        RECT 150.750 104.250 213.750 105.000 ;
        RECT 228.750 104.250 339.750 105.000 ;
        RECT 150.750 103.500 212.250 104.250 ;
        RECT 227.250 103.500 339.000 104.250 ;
        RECT 150.000 102.750 210.750 103.500 ;
        RECT 225.750 102.750 337.500 103.500 ;
        RECT 149.250 102.000 209.250 102.750 ;
        RECT 225.000 102.000 336.750 102.750 ;
        RECT 149.250 101.250 208.500 102.000 ;
        RECT 223.500 101.250 336.000 102.000 ;
        RECT 148.500 100.500 207.000 101.250 ;
        RECT 222.000 100.500 334.500 101.250 ;
        RECT 147.750 99.750 205.500 100.500 ;
        RECT 220.500 99.750 333.750 100.500 ;
        RECT 147.750 99.000 204.750 99.750 ;
        RECT 219.750 99.000 332.250 99.750 ;
        RECT 147.000 98.250 203.250 99.000 ;
        RECT 218.250 98.250 331.500 99.000 ;
        RECT 147.000 97.500 201.750 98.250 ;
        RECT 216.750 97.500 330.000 98.250 ;
        RECT 146.250 96.750 201.000 97.500 ;
        RECT 215.250 96.750 329.250 97.500 ;
        RECT 145.500 96.000 199.500 96.750 ;
        RECT 214.500 96.000 327.750 96.750 ;
        RECT 145.500 95.250 198.000 96.000 ;
        RECT 213.000 95.250 326.250 96.000 ;
        RECT 144.750 94.500 197.250 95.250 ;
        RECT 212.250 94.500 325.500 95.250 ;
        RECT 144.000 93.750 195.750 94.500 ;
        RECT 210.750 93.750 324.000 94.500 ;
        RECT 144.000 93.000 195.000 93.750 ;
        RECT 209.250 93.000 323.250 93.750 ;
        RECT 143.250 92.250 193.500 93.000 ;
        RECT 208.500 92.250 321.750 93.000 ;
        RECT 143.250 91.500 192.000 92.250 ;
        RECT 207.000 91.500 321.000 92.250 ;
        RECT 142.500 90.750 191.250 91.500 ;
        RECT 206.250 90.750 319.500 91.500 ;
        RECT 141.750 90.000 189.750 90.750 ;
        RECT 204.750 90.000 318.750 90.750 ;
        RECT 141.750 89.250 189.000 90.000 ;
        RECT 203.250 89.250 317.250 90.000 ;
        RECT 141.000 88.500 187.500 89.250 ;
        RECT 202.500 88.500 315.750 89.250 ;
        RECT 141.000 87.750 186.000 88.500 ;
        RECT 201.000 87.750 315.000 88.500 ;
        RECT 140.250 87.000 185.250 87.750 ;
        RECT 200.250 87.000 313.500 87.750 ;
        RECT 139.500 86.250 183.750 87.000 ;
        RECT 198.750 86.250 312.000 87.000 ;
        RECT 139.500 85.500 183.000 86.250 ;
        RECT 198.000 85.500 311.250 86.250 ;
        RECT 138.750 84.750 181.500 85.500 ;
        RECT 196.500 84.750 309.750 85.500 ;
        RECT 138.000 84.000 180.750 84.750 ;
        RECT 195.750 84.000 308.250 84.750 ;
        RECT 138.000 83.250 179.250 84.000 ;
        RECT 194.250 83.250 307.500 84.000 ;
        RECT 137.250 82.500 178.500 83.250 ;
        RECT 193.500 82.500 306.000 83.250 ;
        RECT 137.250 81.750 177.000 82.500 ;
        RECT 192.000 81.750 304.500 82.500 ;
        RECT 136.500 81.000 176.250 81.750 ;
        RECT 191.250 81.000 303.750 81.750 ;
        RECT 135.750 80.250 174.750 81.000 ;
        RECT 189.750 80.250 302.250 81.000 ;
        RECT 135.750 79.500 174.000 80.250 ;
        RECT 189.000 79.500 300.750 80.250 ;
        RECT 135.000 78.750 172.500 79.500 ;
        RECT 187.500 78.750 300.000 79.500 ;
        RECT 135.000 78.000 171.750 78.750 ;
        RECT 186.750 78.000 298.500 78.750 ;
        RECT 134.250 77.250 171.000 78.000 ;
        RECT 185.250 77.250 297.000 78.000 ;
        RECT 134.250 76.500 169.500 77.250 ;
        RECT 184.500 76.500 296.250 77.250 ;
        RECT 133.500 75.750 168.750 76.500 ;
        RECT 183.000 75.750 294.750 76.500 ;
        RECT 132.750 75.000 167.250 75.750 ;
        RECT 182.250 75.000 293.250 75.750 ;
        RECT 132.750 74.250 166.500 75.000 ;
        RECT 180.750 74.250 292.500 75.000 ;
        RECT 132.000 73.500 165.000 74.250 ;
        RECT 180.000 73.500 291.000 74.250 ;
        RECT 132.000 72.750 164.250 73.500 ;
        RECT 178.500 72.750 289.500 73.500 ;
        RECT 131.250 72.000 163.500 72.750 ;
        RECT 177.750 72.000 288.750 72.750 ;
        RECT 130.500 71.250 162.000 72.000 ;
        RECT 176.250 71.250 287.250 72.000 ;
        RECT 130.500 70.500 161.250 71.250 ;
        RECT 175.500 70.500 285.750 71.250 ;
        RECT 129.750 69.750 159.750 70.500 ;
        RECT 174.000 69.750 285.000 70.500 ;
        RECT 129.750 69.000 159.000 69.750 ;
        RECT 173.250 69.000 283.500 69.750 ;
        RECT 129.000 68.250 158.250 69.000 ;
        RECT 171.750 68.250 282.000 69.000 ;
        RECT 129.000 67.500 156.750 68.250 ;
        RECT 171.000 67.500 281.250 68.250 ;
        RECT 128.250 66.750 156.000 67.500 ;
        RECT 169.500 66.750 279.750 67.500 ;
        RECT 128.250 66.000 155.250 66.750 ;
        RECT 168.750 66.000 278.250 66.750 ;
        RECT 127.500 65.250 153.750 66.000 ;
        RECT 167.250 65.250 277.500 66.000 ;
        RECT 127.500 64.500 153.000 65.250 ;
        RECT 166.500 64.500 276.000 65.250 ;
        RECT 126.750 63.750 152.250 64.500 ;
        RECT 165.000 63.750 274.500 64.500 ;
        RECT 126.000 63.000 150.750 63.750 ;
        RECT 164.250 63.000 273.750 63.750 ;
        RECT 126.000 62.250 150.000 63.000 ;
        RECT 162.750 62.250 272.250 63.000 ;
        RECT 125.250 61.500 149.250 62.250 ;
        RECT 162.000 61.500 270.750 62.250 ;
        RECT 125.250 60.750 148.500 61.500 ;
        RECT 160.500 60.750 270.000 61.500 ;
        RECT 124.500 60.000 147.000 60.750 ;
        RECT 159.750 60.000 268.500 60.750 ;
        RECT 124.500 59.250 146.250 60.000 ;
        RECT 158.250 59.250 267.750 60.000 ;
        RECT 123.750 58.500 145.500 59.250 ;
        RECT 157.500 58.500 266.250 59.250 ;
        RECT 123.750 57.750 144.000 58.500 ;
        RECT 156.750 57.750 264.750 58.500 ;
        RECT 123.000 57.000 143.250 57.750 ;
        RECT 155.250 57.000 263.250 57.750 ;
        RECT 123.000 56.250 142.500 57.000 ;
        RECT 154.500 56.250 261.750 57.000 ;
        RECT 122.250 55.500 141.750 56.250 ;
        RECT 153.000 55.500 259.500 56.250 ;
        RECT 122.250 54.750 140.250 55.500 ;
        RECT 152.250 54.750 258.000 55.500 ;
        RECT 121.500 54.000 139.500 54.750 ;
        RECT 150.750 54.000 255.750 54.750 ;
        RECT 121.500 53.250 138.750 54.000 ;
        RECT 150.000 53.250 254.250 54.000 ;
        RECT 121.500 52.500 138.000 53.250 ;
        RECT 149.250 52.500 252.000 53.250 ;
        RECT 120.750 51.750 136.500 52.500 ;
        RECT 147.750 51.750 249.750 52.500 ;
        RECT 120.750 51.000 135.750 51.750 ;
        RECT 147.000 51.000 248.250 51.750 ;
        RECT 120.000 50.250 135.000 51.000 ;
        RECT 145.500 50.250 246.000 51.000 ;
        RECT 262.500 50.250 264.000 51.000 ;
        RECT 120.000 49.500 134.250 50.250 ;
        RECT 144.750 49.500 244.500 50.250 ;
        RECT 260.250 49.500 263.250 50.250 ;
        RECT 119.250 48.750 132.750 49.500 ;
        RECT 143.250 48.750 242.250 49.500 ;
        RECT 258.750 48.750 262.500 49.500 ;
        RECT 119.250 48.000 132.000 48.750 ;
        RECT 142.500 48.000 240.750 48.750 ;
        RECT 256.500 48.000 261.750 48.750 ;
        RECT 119.250 47.250 131.250 48.000 ;
        RECT 141.750 47.250 238.500 48.000 ;
        RECT 254.250 47.250 261.000 48.000 ;
        RECT 118.500 46.500 129.750 47.250 ;
        RECT 140.250 46.500 237.000 47.250 ;
        RECT 252.750 46.500 260.250 47.250 ;
        RECT 118.500 45.750 129.000 46.500 ;
        RECT 139.500 45.750 234.750 46.500 ;
        RECT 250.500 45.750 259.500 46.500 ;
        RECT 117.750 45.000 128.250 45.750 ;
        RECT 138.750 45.000 233.250 45.750 ;
        RECT 248.250 45.000 258.750 45.750 ;
        RECT 117.750 44.250 127.500 45.000 ;
        RECT 137.250 44.250 231.000 45.000 ;
        RECT 246.750 44.250 258.000 45.000 ;
        RECT 117.750 43.500 126.000 44.250 ;
        RECT 136.500 43.500 229.500 44.250 ;
        RECT 244.500 43.500 256.500 44.250 ;
        RECT 117.000 42.750 125.250 43.500 ;
        RECT 135.000 42.750 227.250 43.500 ;
        RECT 242.250 42.750 255.750 43.500 ;
        RECT 117.000 42.000 124.500 42.750 ;
        RECT 134.250 42.000 225.000 42.750 ;
        RECT 240.000 42.000 255.000 42.750 ;
        RECT 116.250 41.250 123.000 42.000 ;
        RECT 133.500 41.250 223.500 42.000 ;
        RECT 238.500 41.250 254.250 42.000 ;
        RECT 116.250 40.500 122.250 41.250 ;
        RECT 132.000 40.500 221.250 41.250 ;
        RECT 236.250 40.500 253.500 41.250 ;
        RECT 116.250 39.750 121.500 40.500 ;
        RECT 131.250 39.750 219.750 40.500 ;
        RECT 234.000 39.750 252.750 40.500 ;
        RECT 115.500 39.000 120.000 39.750 ;
        RECT 130.500 39.000 217.500 39.750 ;
        RECT 232.500 39.000 252.000 39.750 ;
        RECT 115.500 38.250 119.250 39.000 ;
        RECT 129.000 38.250 216.000 39.000 ;
        RECT 230.250 38.250 251.250 39.000 ;
        RECT 115.500 37.500 118.500 38.250 ;
        RECT 128.250 37.500 213.750 38.250 ;
        RECT 228.000 37.500 250.500 38.250 ;
        RECT 114.750 36.750 117.000 37.500 ;
        RECT 127.500 36.750 212.250 37.500 ;
        RECT 226.500 36.750 249.750 37.500 ;
        RECT 114.750 36.000 116.250 36.750 ;
        RECT 126.000 36.000 210.000 36.750 ;
        RECT 224.250 36.000 248.250 36.750 ;
        RECT 114.000 35.250 115.500 36.000 ;
        RECT 125.250 35.250 155.250 36.000 ;
        RECT 222.000 35.250 247.500 36.000 ;
        RECT 124.500 34.500 150.000 35.250 ;
        RECT 220.500 34.500 246.750 35.250 ;
        RECT 123.000 33.750 147.000 34.500 ;
        RECT 218.250 33.750 246.000 34.500 ;
        RECT 122.250 33.000 144.000 33.750 ;
        RECT 216.000 33.000 245.250 33.750 ;
        RECT 121.500 32.250 142.500 33.000 ;
        RECT 214.500 32.250 244.500 33.000 ;
        RECT 120.750 31.500 140.250 32.250 ;
        RECT 212.250 31.500 243.750 32.250 ;
        RECT 120.000 30.750 138.750 31.500 ;
        RECT 188.250 30.750 242.250 31.500 ;
        RECT 118.500 30.000 137.250 30.750 ;
        RECT 185.250 30.000 241.500 30.750 ;
        RECT 117.750 29.250 135.000 30.000 ;
        RECT 183.000 29.250 240.750 30.000 ;
        RECT 117.000 28.500 134.250 29.250 ;
        RECT 180.000 28.500 239.250 29.250 ;
        RECT 116.250 27.750 132.750 28.500 ;
        RECT 176.250 27.750 238.500 28.500 ;
        RECT 115.500 27.000 131.250 27.750 ;
        RECT 171.750 27.000 237.750 27.750 ;
        RECT 114.750 26.250 129.750 27.000 ;
        RECT 165.750 26.250 237.000 27.000 ;
        RECT 114.000 25.500 129.000 26.250 ;
        RECT 136.500 25.500 146.250 26.250 ;
        RECT 155.250 25.500 235.500 26.250 ;
        RECT 113.250 24.750 127.500 25.500 ;
        RECT 135.750 24.750 234.750 25.500 ;
        RECT 112.500 24.000 126.750 24.750 ;
        RECT 135.000 24.000 233.250 24.750 ;
        RECT 111.750 23.250 125.250 24.000 ;
        RECT 133.500 23.250 232.500 24.000 ;
        RECT 111.000 22.500 124.500 23.250 ;
        RECT 132.750 22.500 231.000 23.250 ;
        RECT 110.250 21.750 123.000 22.500 ;
        RECT 132.000 21.750 230.250 22.500 ;
        RECT 110.250 21.000 122.250 21.750 ;
        RECT 131.250 21.000 228.750 21.750 ;
        RECT 109.500 20.250 121.500 21.000 ;
        RECT 130.500 20.250 228.000 21.000 ;
        RECT 108.750 19.500 120.000 20.250 ;
        RECT 129.000 19.500 226.500 20.250 ;
        RECT 108.750 18.750 119.250 19.500 ;
        RECT 128.250 18.750 225.000 19.500 ;
        RECT 108.000 18.000 118.500 18.750 ;
        RECT 127.500 18.000 224.250 18.750 ;
        RECT 107.250 17.250 117.000 18.000 ;
        RECT 126.750 17.250 222.750 18.000 ;
        RECT 107.250 16.500 116.250 17.250 ;
        RECT 125.250 16.500 221.250 17.250 ;
        RECT 106.500 15.750 115.500 16.500 ;
        RECT 124.500 15.750 219.750 16.500 ;
        RECT 106.500 15.000 114.000 15.750 ;
        RECT 123.750 15.000 218.250 15.750 ;
        RECT 105.750 14.250 113.250 15.000 ;
        RECT 123.000 14.250 216.750 15.000 ;
        RECT 105.750 13.500 111.750 14.250 ;
        RECT 121.500 13.500 215.250 14.250 ;
        RECT 105.000 12.750 111.000 13.500 ;
        RECT 120.750 12.750 213.750 13.500 ;
        RECT 105.000 12.000 109.500 12.750 ;
        RECT 120.000 12.000 212.250 12.750 ;
        RECT 104.250 11.250 108.750 12.000 ;
        RECT 119.250 11.250 210.000 12.000 ;
        RECT 104.250 10.500 107.250 11.250 ;
        RECT 118.500 10.500 208.500 11.250 ;
        RECT 103.500 9.750 105.750 10.500 ;
        RECT 117.000 9.750 206.250 10.500 ;
        RECT 103.500 9.000 105.000 9.750 ;
        RECT 116.250 9.000 204.750 9.750 ;
        RECT 115.500 8.250 202.500 9.000 ;
        RECT 114.750 7.500 200.250 8.250 ;
        RECT 113.250 6.750 198.000 7.500 ;
        RECT 112.500 6.000 195.750 6.750 ;
        RECT 111.750 5.250 192.750 6.000 ;
        RECT 114.750 4.500 190.500 5.250 ;
        RECT 119.250 3.750 187.500 4.500 ;
        RECT 124.500 3.000 183.750 3.750 ;
        RECT 129.000 2.250 180.750 3.000 ;
        RECT 135.000 1.500 176.250 2.250 ;
        RECT 141.000 0.750 171.000 1.500 ;
        RECT 151.500 0.000 160.500 0.750 ;
  END
END avali_logo
END LIBRARY

